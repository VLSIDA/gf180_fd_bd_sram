* Subcircuit definition of cell ICV_19
.SUBCKT ICV_19
** N=6 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
