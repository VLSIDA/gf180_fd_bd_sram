* Subcircuit definition of cell mux821
.SUBCKT mux821 1 2 3 4 5 6 7 8 9 13 14 15 16 17 18 19 20 21 22 23
+ 24 25 26 27 28 29 30 31 32 33 42 43 44 45 46 47 48
** N=86 EP=37 IP=165 FDC=48
*.SEEDPROM
M0 13 42 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=1510 $Y=2370 $D=2
M1 16 43 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=3750 $Y=2370 $D=2
M2 19 44 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=7705 $Y=2370 $D=2
M3 22 45 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=9945 $Y=2370 $D=2
M4 25 46 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=13895 $Y=2370 $D=2
M5 28 47 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=16135 $Y=2370 $D=2
M6 31 48 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=20090 $Y=2370 $D=2
M7 2 9 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=22330 $Y=2370 $D=2
X9 5 3 7 8 pfet_05v0_I01 $T=23310 51440 1 0 $X=22270 $Y=44010
X10 5 6 2 8 pfet_05v0_I01 $T=23320 43505 1 0 $X=22280 $Y=36075
X12 3 4 2 8 pmos_1p2$$46889004 $T=23475 15755 1 0 $X=22045 $Y=8245
X13 3 4 9 1 nmos_1p2$$47119404 $T=23475 25030 1 0 $X=22330 $Y=17545
X14 5 6 9 1 nmos_1p2$$47119404 $T=23475 35050 1 0 $X=22330 $Y=27565
X15 1 13 15 4 14 6 42 7 8 ypass_gate $T=3490 455 1 180 $X=-1160 $Y=0
X16 1 16 18 4 17 6 43 7 8 ypass_gate $T=3490 455 0 0 $X=2385 $Y=0
X17 1 19 21 4 20 6 44 7 8 ypass_gate $T=9685 455 1 180 $X=5035 $Y=0
X18 1 22 24 4 23 6 45 7 8 ypass_gate $T=9685 455 0 0 $X=8580 $Y=0
X19 1 25 27 4 26 6 46 7 8 ypass_gate $T=15875 455 1 180 $X=11225 $Y=0
X20 1 28 30 4 29 6 47 7 8 ypass_gate $T=15875 455 0 0 $X=14770 $Y=0
X21 1 31 33 4 32 6 48 7 8 ypass_gate $T=22070 455 1 180 $X=17420 $Y=0
.ENDS
