* Subcircuit definition of cell ICV_13
.SUBCKT ICV_13 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=26 EP=17 IP=30 FDC=16
*.SEEDPROM
X0 1 1 3 4 5 6 7 8 9 10 ICV_6 $T=-6000 0 0 0 $X=-9340 $Y=-340
X1 1 1 11 12 13 14 15 16 17 18 ICV_6 $T=0 0 0 0 $X=-3340 $Y=-340
.ENDS
