* Subcircuit definition of cell nfet_05v0_I12
.SUBCKT nfet_05v0_I12
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
