* Subcircuit definition of cell pmos_1p2$$46898220
.SUBCKT pmos_1p2$$46898220
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
