* Subcircuit definition of cell pfet_05v0_I14
.SUBCKT pfet_05v0_I14
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
