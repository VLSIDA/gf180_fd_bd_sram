* Subcircuit definition of cell xpredec1
.SUBCKT xpredec1 vss men vdd clk A[2] A[1] A[0] x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0]
** N=91 EP=15 IP=199 FDC=108
M0 77 18 51 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=1700 $Y=2310 $D=2
M1 76 19 77 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=2820 $Y=2310 $D=2
M2 vss 20 76 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=3940 $Y=2310 $D=2
M3 vss 51 x[7] vss nfet_05v0 L=6e-07 W=1.362e-05 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=1700 $Y=48000 $D=2
M4 78 21 vss vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=5060 $Y=2310 $D=2
M5 79 19 78 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=6180 $Y=2310 $D=2
M6 54 18 79 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=7300 $Y=2310 $D=2
M7 x[6] 54 vss vss nfet_05v0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=5060 $Y=48000 $D=2
M8 81 18 57 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=9870 $Y=2310 $D=2
M9 80 22 81 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=10990 $Y=2310 $D=2
M10 vss 20 80 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12110 $Y=2310 $D=2
M11 vss 57 x[5] vss nfet_05v0 L=6e-07 W=1.362e-05 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=9870 $Y=48000 $D=2
M12 82 21 vss vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=13230 $Y=2310 $D=2
M13 83 22 82 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=14350 $Y=2310 $D=2
M14 60 18 83 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=15470 $Y=2310 $D=2
M15 x[4] 60 vss vss nfet_05v0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=13230 $Y=48000 $D=2
M16 85 23 63 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=18035 $Y=2310 $D=2
M17 84 19 85 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=19155 $Y=2310 $D=2
M18 vss 20 84 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=20275 $Y=2310 $D=2
M19 vss 63 x[3] vss nfet_05v0 L=6e-07 W=1.362e-05 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=18035 $Y=48000 $D=2
M20 86 21 vss vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=21395 $Y=2310 $D=2
M21 87 19 86 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=22515 $Y=2310 $D=2
M22 66 23 87 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=23635 $Y=2310 $D=2
M23 x[2] 66 vss vss nfet_05v0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=21395 $Y=48000 $D=2
M24 89 23 69 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=26205 $Y=2310 $D=2
M25 88 22 89 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=27325 $Y=2310 $D=2
M26 vss 20 88 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=28445 $Y=2310 $D=2
M27 vss 69 x[1] vss nfet_05v0 L=6e-07 W=1.362e-05 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=26205 $Y=48000 $D=2
M28 90 21 vss vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=29565 $Y=2310 $D=2
M29 91 22 90 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=30685 $Y=2310 $D=2
M30 72 23 91 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=31805 $Y=2310 $D=2
M31 x[0] 72 vss vss nfet_05v0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=29565 $Y=48000 $D=2
M32 17 men vss vss nfet_05v0 L=6e-07 W=1.91e-06 AD=4.966e-13 AS=8.404e-13 PD=2.43e-06 PS=4.7e-06 NRD=0.136126 NRS=0.230366 m=1 nf=1 $X=37165 $Y=51200 $D=2
M33 vss clk 17 vss nfet_05v0 L=6e-07 W=1.91e-06 AD=8.404e-13 AS=4.966e-13 PD=4.7e-06 PS=2.43e-06 NRD=0.230366 NRS=0.136126 m=1 nf=1 $X=38285 $Y=51200 $D=2
M34 vss 17 16 vss nfet_05v0 L=6e-07 W=1.36e-06 AD=5.984e-13 AS=5.984e-13 PD=3.6e-06 PS=3.6e-06 NRD=0.323529 NRS=0.323529 m=1 nf=1 $X=45140 $Y=51180 $D=2
M35 vdd 18 51 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=1700 $Y=21650 $D=8
M36 51 19 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=2820 $Y=21650 $D=8
M37 vdd 20 51 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=3940 $Y=21650 $D=8
M38 vdd 51 x[7] vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=1700 $Y=35260 $D=8
M39 54 21 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=5060 $Y=21650 $D=8
M40 vdd 19 54 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=6180 $Y=21650 $D=8
M41 54 18 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=7300 $Y=21650 $D=8
M42 x[6] 54 vdd vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=5060 $Y=35260 $D=8
M43 vdd 18 57 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=9870 $Y=21650 $D=8
M44 57 22 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=10990 $Y=21650 $D=8
M45 vdd 20 57 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12110 $Y=21650 $D=8
M46 vdd 57 x[5] vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=9870 $Y=35260 $D=8
M47 60 21 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=13230 $Y=21650 $D=8
M48 vdd 22 60 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=14350 $Y=21650 $D=8
M49 60 18 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=15470 $Y=21650 $D=8
M50 x[4] 60 vdd vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=13230 $Y=35260 $D=8
M51 vdd 23 63 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=18035 $Y=21650 $D=8
M52 63 19 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=19155 $Y=21650 $D=8
M53 vdd 20 63 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=20275 $Y=21650 $D=8
M54 vdd 63 x[3] vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=18035 $Y=35260 $D=8
M55 66 21 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=21395 $Y=21650 $D=8
M56 vdd 19 66 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=22515 $Y=21650 $D=8
M57 66 23 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=23635 $Y=21650 $D=8
M58 x[2] 66 vdd vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=21395 $Y=35260 $D=8
M59 vdd 23 69 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=26205 $Y=21650 $D=8
M60 69 22 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=27325 $Y=21650 $D=8
M61 vdd 20 69 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=28445 $Y=21650 $D=8
M62 vdd 69 x[1] vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=26205 $Y=35260 $D=8
M63 72 21 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=29565 $Y=21650 $D=8
M64 vdd 22 72 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=30685 $Y=21650 $D=8
M65 72 23 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=31805 $Y=21650 $D=8
M66 x[0] 72 vdd vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=29565 $Y=35260 $D=8
M67 74 men vdd vdd pfet_05v0 L=6e-07 W=2.275e-06 AD=5.915e-13 AS=1.35362e-12 PD=2.795e-06 PS=5.74e-06 NRD=0.114286 NRS=0.261538 m=1 nf=1 $X=37165 $Y=47525 $D=8
M68 17 clk 74 vdd pfet_05v0 L=6e-07 W=2.275e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=38285 $Y=47525 $D=8
M69 75 clk 17 vdd pfet_05v0 L=6e-07 W=2.275e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=39405 $Y=47525 $D=8
M70 vdd men 75 vdd pfet_05v0 L=6e-07 W=2.275e-06 AD=1.35362e-12 AS=5.915e-13 PD=5.74e-06 PS=2.795e-06 NRD=0.261538 NRS=0.114286 m=1 nf=1 $X=40525 $Y=47525 $D=8
X71 vdd 16 17 pmos_1p2$$47109164 $T=44700 47595 0 0 $X=42105 $Y=46910
X83 vss 18 23 vdd A[2] 17 16 xpredec1_bot $T=34205 3160 0 0 $X=33675 $Y=-5
X84 vss 19 22 vdd A[1] 17 16 xpredec1_bot $T=42655 3160 0 0 $X=42125 $Y=-5
X85 vss 20 21 vdd A[0] 17 16 xpredec1_bot $T=51110 3160 0 0 $X=50580 $Y=-5
.ENDS
