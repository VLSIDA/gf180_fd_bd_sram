* Subcircuit definition of cell ICV_3
.SUBCKT ICV_3 1 2 3 4 10 12 14 15
** N=19 EP=8 IP=26 FDC=16
*.SEEDPROM
M0 1 3 16 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=3180 $Y=7970 $D=2
M1 18 3 1 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=3180 $Y=9260 $D=2
M2 3 4 16 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=3630 $Y=6340 $D=2
M3 3 4 18 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=3630 $Y=10710 $D=2
M4 17 3 3 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=4770 $Y=6340 $D=2
M5 19 3 3 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=4770 $Y=10710 $D=2
M6 2 3 17 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=5220 $Y=7970 $D=2
M7 19 3 2 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=5220 $Y=9260 $D=2
X8 3 4 10 12 16 17 ICV_2 $T=0 0 0 0 $X=-340 $Y=-340
X9 3 4 18 19 14 15 ICV_2 $T=0 9000 0 0 $X=-340 $Y=8660
.ENDS
