* Subcircuit definition of cell ICV_12
.SUBCKT ICV_12
** N=27 EP=0 IP=32 FDC=0
.ENDS
