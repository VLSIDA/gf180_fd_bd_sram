* Subcircuit definition of cell gf180mcu_fd_ip_sram__sram128x8m8wm1
.SUBCKT gf180mcu_fd_ip_sram__sram128x8m8wm1 A[6] A[5] A[4] A[3] A[2] A[1] A[0]
+ CEN CLK D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] GWEN Q[7] Q[6] Q[5] Q[4]
+ Q[3] Q[2] Q[1] Q[0] VDD VSS WEN[7] WEN[6] WEN[5] WEN[4] WEN[3] WEN[2] WEN[1]
+ WEN[0]
** N=5565 EP=36 IP=3508 FDC=9725
M0 4646 VSS 733 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=120390 $Y=176390 $D=2
M1 733 VSS 4648 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=120390 $Y=256100 $D=2
M2 VSS 4645 4646 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=120840 $Y=177840 $D=2
M3 VSS 4647 4648 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=120840 $Y=254470 $D=2
M4 4645 4646 VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=121980 $Y=177840 $D=2
M5 4647 4648 VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=121980 $Y=254470 $D=2
M6 4645 VSS 732 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=122430 $Y=176390 $D=2
M7 732 VSS 4647 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=122430 $Y=256100 $D=2
M8 VSS 4854 4222 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=168355 $Y=180895 $D=2
M9 4854 4826 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=183295 $D=2
M10 VSS 4828 4856 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=213375 $D=2
M11 VSS 4856 4229 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=214655 $D=2
M12 VSS 4858 4230 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=216895 $D=2
M13 4858 4830 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=219295 $D=2
M14 VSS 4832 4860 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=249375 $D=2
M15 VSS 4860 4237 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=168355 $Y=250655 $D=2
M16 4826 4827 VSS VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=198635 $Y=180895 $D=2
M17 VSS 4829 4828 VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=215775 $D=2
M18 4830 4831 VSS VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=216895 $D=2
M19 VSS 4833 4832 VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=198635 $Y=251775 $D=2
M20 2 VDD 1 VSS nfet_05v0 L=6e-07 W=6.59e-06 AD=2.8996e-12 AS=2.8996e-12 PD=1.406e-05 PS=1.406e-05 NRD=0.0667678 NRS=0.0667678 m=1 nf=1 $X=204815 $Y=255000 $D=2
M21 5527 VDD VSS VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=7.32375e-13 AS=2.079e-12 PD=3.615e-06 PS=7.62e-06 NRD=0.0738095 NRS=0.209524 m=1 nf=1 $X=218475 $Y=180950 $D=2
M22 5526 918 5527 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=182015 $D=2
M23 4827 926 5526 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=183135 $D=2
M24 5528 919 4829 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=213535 $D=2
M25 5529 918 5528 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=214655 $D=2
M26 VSS VDD 5529 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=215720 $D=2
M27 5531 VDD VSS VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=216950 $D=2
M28 5530 917 5531 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=218015 $D=2
M29 4831 926 5530 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=219135 $D=2
M30 5532 919 4833 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=249535 $D=2
M31 5533 917 5532 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=250655 $D=2
M32 VSS VDD 5533 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.079e-12 AS=7.32375e-13 PD=7.62e-06 PS=3.615e-06 NRD=0.209524 NRS=0.0738095 m=1 nf=1 $X=218475 $Y=251720 $D=2
M33 VSS 1 787 VSS nfet_05v0 L=6e-07 W=1.36e-06 AD=3.536e-13 AS=5.984e-13 PD=1.88e-06 PS=3.6e-06 NRD=0.191176 NRS=0.323529 m=1 nf=1 $X=233770 $Y=54135 $D=2
M34 787 CLK VSS VSS nfet_05v0 L=6e-07 W=1.36e-06 AD=5.984e-13 AS=3.536e-13 PD=3.6e-06 PS=1.88e-06 NRD=0.323529 NRS=0.191176 m=1 nf=1 $X=234890 $Y=54135 $D=2
M35 616 619 VSS VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=242235 $Y=54135 $D=2
M36 281 865 VSS VSS nfet_05v0 L=1e-06 W=6e-07 AD=2.64e-13 AS=2.64e-13 PD=2.08e-06 PS=2.08e-06 NRD=0.733333 NRS=0.733333 m=1 nf=1 $X=243265 $Y=46010 $D=2
M37 CEN 787 619 VSS nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=245925 $Y=54135 $D=2
M38 250 468 VSS VSS nfet_05v0 L=6e-07 W=4.99e-05 AD=1.47704e-11 AS=1.47704e-11 PD=6.284e-05 PS=6.284e-05 NRD=0.148297 NRS=0.148297 m=1 nf=5 $X=241995 $Y=72320 $D=2
M39 317 281 VSS VSS nfet_05v0 L=6e-07 W=7.5e-07 AD=3.3e-13 AS=3.3e-13 PD=2.38e-06 PS=2.38e-06 NRD=0.586667 NRS=0.586667 m=1 nf=1 $X=246495 $Y=46075 $D=2
M40 354 317 VSS VSS nfet_05v0 L=6e-07 W=3.02e-06 AD=1.3288e-12 AS=1.3288e-12 PD=6.92e-06 PS=6.92e-06 NRD=0.145695 NRS=0.145695 m=1 nf=1 $X=249065 $Y=46070 $D=2
M41 4811 354 VSS VSS nfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=1.34946e-11 PD=2.32e-05 PS=4.655e-05 NRD=0.0114638 NRS=0.0262346 m=1 nf=1 $X=256125 $Y=28435 $D=2
M42 VSS 4855 4238 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=252270 $Y=180895 $D=2
M43 4855 4826 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=183295 $D=2
M44 VSS 4828 4857 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=213375 $D=2
M45 VSS 4857 4245 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=214655 $D=2
M46 VSS 4859 4246 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=216895 $D=2
M47 4859 4830 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=219295 $D=2
M48 VSS 4832 4861 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=249375 $D=2
M49 VSS 4861 4253 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=252270 $Y=250655 $D=2
M50 4812 CLK 4811 VSS nfet_05v0 L=6e-07 W=2.268e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=257245 $Y=28435 $D=2
M51 445 616 4812 VSS nfet_05v0 L=6e-07 W=2.268e-05 AD=1.33812e-11 AS=5.8968e-12 PD=4.654e-05 PS=2.32e-05 NRD=0.0260141 NRS=0.0114638 m=1 nf=1 $X=258365 $Y=28435 $D=2
M52 4813 495 VSS VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=4.7177e-12 AS=1.07963e-11 PD=1.8665e-05 PS=3.748e-05 NRD=0.014329 NRS=0.0327914 m=1 nf=1 $X=262120 $Y=29545 $D=2
M53 468 445 4813 VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=263240 $Y=29545 $D=2
M54 4814 445 468 VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=264360 $Y=29545 $D=2
M55 VSS 495 4814 VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=1.07055e-11 AS=4.7177e-12 PD=3.747e-05 PS=1.8665e-05 NRD=0.0325158 NRS=0.014329 m=1 nf=1 $X=265480 $Y=29545 $D=2
M56 4815 468 VSS VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=1.16905e-12 AS=2.7013e-12 PD=5.055e-06 PS=1.027e-05 NRD=0.0567181 NRS=0.131057 m=1 nf=1 $X=268545 $Y=43150 $D=2
M57 495 607 4815 VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=2.27e-14 AS=-2.27e-14 PD=1e-08 PS=-1e-08 NRD=0.00110132 NRS=-0.00110132 m=1 nf=1 $X=269660 $Y=43150 $D=2
M58 4816 607 495 VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=-2.27e-14 AS=2.27e-14 PD=-1e-08 PS=1e-08 NRD=-0.00110132 NRS=0.00110132 m=1 nf=1 $X=270785 $Y=43150 $D=2
M59 VSS 468 4816 VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=2.7013e-12 AS=1.16905e-12 PD=1.027e-05 PS=5.055e-06 NRD=0.131057 NRS=0.0567181 m=1 nf=1 $X=271900 $Y=43150 $D=2
M60 1 250 VSS VSS nfet_05v0 L=6e-07 W=0.0001474 AD=3.8324e-11 AS=4.09772e-11 PD=0.0001578 PS=0.00017326 NRD=0.705563 NRS=0.75441 m=1 nf=20 $X=253180 $Y=76320 $D=2
M61 4650 VSS 735 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=304270 $Y=176390 $D=2
M62 735 VSS 4652 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=304270 $Y=256100 $D=2
M63 VSS 4649 4650 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=304720 $Y=177840 $D=2
M64 VSS 4651 4652 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=304720 $Y=254470 $D=2
M65 4649 4650 VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=305860 $Y=177840 $D=2
M66 4651 4652 VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=305860 $Y=254470 $D=2
M67 4649 VSS 734 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=306310 $Y=176390 $D=2
M68 734 VSS 4651 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=306310 $Y=256100 $D=2
M69 4838 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=418270 $Y=176390 $D=2
M70 614 VSS 4840 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=193100 $D=2
M71 4842 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=194390 $D=2
M72 614 VSS 4844 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=211100 $D=2
M73 4846 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=212390 $D=2
M74 614 VSS 4848 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=229100 $D=2
M75 4850 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=230390 $D=2
M76 614 861 4852 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=247100 $D=2
M77 4834 861 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=248390 $D=2
M78 614 861 4836 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=418270 $Y=256100 $D=2
M79 VSS VDD 4838 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=177840 $D=2
M80 VSS VDD 4840 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=191470 $D=2
M81 VSS VDD 4842 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=195840 $D=2
M82 VSS VDD 4844 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=209470 $D=2
M83 VSS VDD 4846 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=213840 $D=2
M84 VSS VDD 4848 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=227470 $D=2
M85 VSS VDD 4850 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=231840 $D=2
M86 VSS VDD 4852 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=245470 $D=2
M87 VSS VDD 4834 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=249840 $D=2
M88 VSS VDD 4836 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=254470 $D=2
M89 4839 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=177840 $D=2
M90 4841 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=191470 $D=2
M91 4843 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=195840 $D=2
M92 4845 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=209470 $D=2
M93 4847 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=213840 $D=2
M94 4849 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=227470 $D=2
M95 4851 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=231840 $D=2
M96 4853 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=245470 $D=2
M97 4835 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=249840 $D=2
M98 4837 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=254470 $D=2
M99 606 614 VSS VSS nfet_05v0 L=6e-07 W=2.76e-06 AD=7.176e-13 AS=1.2144e-12 PD=3.8e-06 PS=7.28e-06 NRD=0.376812 NRS=0.637681 m=1 nf=2 $X=418770 $Y=94540 $D=2
M100 607 606 VSS VSS nfet_05v0 L=6e-07 W=1.7e-05 AD=4.42e-12 AS=7.48e-12 PD=1.804e-05 PS=3.576e-05 NRD=0.0611765 NRS=0.103529 m=1 nf=2 $X=418790 $Y=79115 $D=2
M101 613 VDD VSS VSS nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=5.016e-13 PD=2.18e-06 PS=4.04e-06 NRD=0.912281 NRS=1.54386 m=1 nf=2 $X=419015 $Y=110805 $D=2
M102 4839 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=420310 $Y=176390 $D=2
M103 615 VSS 4841 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=193100 $D=2
M104 4843 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=194390 $D=2
M105 615 VSS 4845 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=211100 $D=2
M106 4847 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=212390 $D=2
M107 615 VSS 4849 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=229100 $D=2
M108 4851 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=230390 $D=2
M109 615 861 4853 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=247100 $D=2
M110 4835 861 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=248390 $D=2
M111 615 861 4837 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=420310 $Y=256100 $D=2
M112 VDD 4482 4484 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=179690 $D=8
M113 VDD 4891 4890 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=180970 $D=8
M114 VDD 4899 4898 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=215690 $D=8
M115 VDD 4955 4954 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=216970 $D=8
M116 VDD 4963 4962 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=251690 $D=8
M117 VDD 4498 4500 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=252970 $D=8
M118 4482 4484 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=179690 $D=8
M119 4891 4890 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=180970 $D=8
M120 4899 4898 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=215690 $D=8
M121 4955 4954 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=216970 $D=8
M122 4963 4962 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=251690 $D=8
M123 4498 4500 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=252970 $D=8
M124 4699 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=13620 $Y=160970 $D=8
M125 4700 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=13620 $Y=164845 $D=8
M126 4862 4664 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=13835 $Y=112830 $D=8
M127 VDD 4478 4480 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=179690 $D=8
M128 VDD 4893 4892 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=180970 $D=8
M129 VDD 4901 4900 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=215690 $D=8
M130 VDD 4957 4956 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=216970 $D=8
M131 VDD 4965 4964 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=251690 $D=8
M132 VDD 4494 4496 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=252970 $D=8
M133 4478 4480 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=179690 $D=8
M134 4893 4892 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=180970 $D=8
M135 4901 4900 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=215690 $D=8
M136 4957 4956 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=216970 $D=8
M137 4965 4964 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=251690 $D=8
M138 4494 4496 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=252970 $D=8
M139 4863 4663 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=16365 $Y=112830 $D=8
M140 4702 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=16720 $Y=160970 $D=8
M141 4701 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=16720 $Y=164845 $D=8
M142 VDD 4474 4476 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=179690 $D=8
M143 VDD 4895 4894 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=180970 $D=8
M144 VDD 4903 4902 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=215690 $D=8
M145 VDD 4959 4958 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=216970 $D=8
M146 VDD 4967 4966 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=251690 $D=8
M147 VDD 4490 4492 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=252970 $D=8
M148 4474 4476 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=179690 $D=8
M149 4895 4894 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=180970 $D=8
M150 4903 4902 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=215690 $D=8
M151 4959 4958 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=216970 $D=8
M152 4967 4966 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=251690 $D=8
M153 4490 4492 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=252970 $D=8
M154 4703 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=19815 $Y=160970 $D=8
M155 4704 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=19815 $Y=164845 $D=8
M156 4864 4662 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=20030 $Y=112830 $D=8
M157 VDD 4470 4472 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=179690 $D=8
M158 VDD 4897 4896 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=180970 $D=8
M159 VDD 4905 4904 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=215690 $D=8
M160 VDD 4961 4960 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=216970 $D=8
M161 VDD 4969 4968 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=251690 $D=8
M162 VDD 4486 4488 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=252970 $D=8
M163 4470 4472 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=179690 $D=8
M164 4897 4896 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=180970 $D=8
M165 4905 4904 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=215690 $D=8
M166 4961 4960 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=216970 $D=8
M167 4969 4968 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=251690 $D=8
M168 4486 4488 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=252970 $D=8
M169 4865 4661 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=22560 $Y=112830 $D=8
M170 4706 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=22915 $Y=160970 $D=8
M171 4705 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=22915 $Y=164845 $D=8
M172 VDD 4266 4268 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=179690 $D=8
M173 VDD 4907 4906 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=180970 $D=8
M174 VDD 4915 4914 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=215690 $D=8
M175 VDD 4971 4970 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=216970 $D=8
M176 VDD 4979 4978 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=251690 $D=8
M177 VDD 4338 4340 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=252970 $D=8
M178 4266 4268 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=179690 $D=8
M179 4907 4906 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=180970 $D=8
M180 4915 4914 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=215690 $D=8
M181 4971 4970 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=216970 $D=8
M182 4979 4978 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=251690 $D=8
M183 4338 4340 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=252970 $D=8
M184 4707 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=26005 $Y=160970 $D=8
M185 4708 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=26005 $Y=164845 $D=8
M186 4866 4660 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=26220 $Y=112830 $D=8
M187 VDD 4262 4264 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=179690 $D=8
M188 VDD 4909 4908 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=180970 $D=8
M189 VDD 4917 4916 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=215690 $D=8
M190 VDD 4973 4972 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=216970 $D=8
M191 VDD 4981 4980 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=251690 $D=8
M192 VDD 4334 4336 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=252970 $D=8
M193 4262 4264 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=179690 $D=8
M194 4909 4908 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=180970 $D=8
M195 4917 4916 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=215690 $D=8
M196 4973 4972 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=216970 $D=8
M197 4981 4980 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=251690 $D=8
M198 4334 4336 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=252970 $D=8
M199 4867 4659 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=28750 $Y=112830 $D=8
M200 4710 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=29105 $Y=160970 $D=8
M201 4709 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=29105 $Y=164845 $D=8
M202 VDD 4274 4276 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=179690 $D=8
M203 VDD 4911 4910 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=180970 $D=8
M204 VDD 4919 4918 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=215690 $D=8
M205 VDD 4975 4974 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=216970 $D=8
M206 VDD 4983 4982 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=251690 $D=8
M207 VDD 4330 4332 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=252970 $D=8
M208 4274 4276 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=179690 $D=8
M209 4911 4910 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=180970 $D=8
M210 4919 4918 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=215690 $D=8
M211 4975 4974 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=216970 $D=8
M212 4983 4982 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=251690 $D=8
M213 4330 4332 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=252970 $D=8
M214 4711 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=32200 $Y=160970 $D=8
M215 4712 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=32200 $Y=164845 $D=8
M216 4868 4658 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=32415 $Y=112830 $D=8
M217 VDD 4270 4272 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=179690 $D=8
M218 VDD 4913 4912 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=180970 $D=8
M219 VDD 4921 4920 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=215690 $D=8
M220 VDD 4977 4976 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=216970 $D=8
M221 VDD 4985 4984 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=251690 $D=8
M222 VDD 4326 4328 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=252970 $D=8
M223 4270 4272 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=179690 $D=8
M224 4913 4912 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=180970 $D=8
M225 4921 4920 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=215690 $D=8
M226 4977 4976 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=216970 $D=8
M227 4985 4984 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=251690 $D=8
M228 4326 4328 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=252970 $D=8
M229 4818 4657 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=34945 $Y=112830 $D=8
M230 938 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=35120 $Y=160970 $D=8
M231 939 4218 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=35120 $Y=164845 $D=8
M232 950 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=38575 $Y=160970 $D=8
M233 951 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=38575 $Y=164845 $D=8
M234 VDD 4514 4516 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=179690 $D=8
M235 VDD 4928 4929 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=180970 $D=8
M236 VDD 4936 4937 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=215690 $D=8
M237 VDD 4992 4993 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=216970 $D=8
M238 VDD 5000 5001 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=251690 $D=8
M239 VDD 4530 4532 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=252970 $D=8
M240 4822 4664 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=38620 $Y=112830 $D=8
M241 4514 4516 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=179690 $D=8
M242 4928 4929 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=180970 $D=8
M243 4936 4937 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=215690 $D=8
M244 4992 4993 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=216970 $D=8
M245 5000 5001 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=251690 $D=8
M246 4530 4532 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=252970 $D=8
M247 5408 4663 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=41145 $Y=112830 $D=8
M248 4791 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=41500 $Y=160970 $D=8
M249 4792 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=41500 $Y=164845 $D=8
M250 VDD 4510 4512 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=179690 $D=8
M251 VDD 4926 4927 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=180970 $D=8
M252 VDD 4934 4935 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=215690 $D=8
M253 VDD 4990 4991 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=216970 $D=8
M254 VDD 4998 4999 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=251690 $D=8
M255 VDD 4526 4528 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=252970 $D=8
M256 4510 4512 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=179690 $D=8
M257 4926 4927 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=180970 $D=8
M258 4934 4935 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=215690 $D=8
M259 4990 4991 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=216970 $D=8
M260 4998 4999 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=251690 $D=8
M261 4526 4528 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=252970 $D=8
M262 4790 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=44595 $Y=160970 $D=8
M263 4789 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=44595 $Y=164845 $D=8
M264 VDD 4506 4508 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=179690 $D=8
M265 VDD 4924 4925 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=180970 $D=8
M266 VDD 4932 4933 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=215690 $D=8
M267 VDD 4988 4989 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=216970 $D=8
M268 VDD 4996 4997 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=251690 $D=8
M269 VDD 4522 4524 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=252970 $D=8
M270 5407 4662 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=44810 $Y=112830 $D=8
M271 4506 4508 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=179690 $D=8
M272 4924 4925 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=180970 $D=8
M273 4932 4933 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=215690 $D=8
M274 4988 4989 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=216970 $D=8
M275 4996 4997 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=251690 $D=8
M276 4522 4524 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=252970 $D=8
M277 5406 4661 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=47340 $Y=112830 $D=8
M278 4787 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=47695 $Y=160970 $D=8
M279 4788 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=47695 $Y=164845 $D=8
M280 VDD 4502 4504 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=179690 $D=8
M281 VDD 4922 4923 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=180970 $D=8
M282 VDD 4930 4931 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=215690 $D=8
M283 VDD 4986 4987 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=216970 $D=8
M284 VDD 4994 4995 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=251690 $D=8
M285 VDD 4518 4520 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=252970 $D=8
M286 4502 4504 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=179690 $D=8
M287 4922 4923 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=180970 $D=8
M288 4930 4931 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=215690 $D=8
M289 4986 4987 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=216970 $D=8
M290 4994 4995 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=251690 $D=8
M291 4518 4520 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=252970 $D=8
M292 VDD 4354 4356 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=179690 $D=8
M293 VDD 4944 4945 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=180970 $D=8
M294 VDD 4952 4953 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=215690 $D=8
M295 VDD 5008 5009 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=216970 $D=8
M296 VDD 5016 5017 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=251690 $D=8
M297 VDD 4370 4372 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=252970 $D=8
M298 4762 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=50785 $Y=160970 $D=8
M299 4761 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=50785 $Y=164845 $D=8
M300 5405 4660 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=51000 $Y=112830 $D=8
M301 4354 4356 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=179690 $D=8
M302 4944 4945 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=180970 $D=8
M303 4952 4953 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=215690 $D=8
M304 5008 5009 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=216970 $D=8
M305 5016 5017 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=251690 $D=8
M306 4370 4372 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=252970 $D=8
M307 5404 4659 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=53530 $Y=112830 $D=8
M308 VDD 4350 4352 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=179690 $D=8
M309 VDD 4942 4943 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=180970 $D=8
M310 VDD 4950 4951 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=215690 $D=8
M311 VDD 5006 5007 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=216970 $D=8
M312 VDD 5014 5015 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=251690 $D=8
M313 VDD 4366 4368 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=252970 $D=8
M314 4759 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=53885 $Y=160970 $D=8
M315 4760 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=53885 $Y=164845 $D=8
M316 4350 4352 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=179690 $D=8
M317 4942 4943 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=180970 $D=8
M318 4950 4951 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=215690 $D=8
M319 5006 5007 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=216970 $D=8
M320 5014 5015 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=251690 $D=8
M321 4366 4368 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=252970 $D=8
M322 VDD 4346 4348 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=179690 $D=8
M323 VDD 4940 4941 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=180970 $D=8
M324 VDD 4948 4949 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=215690 $D=8
M325 VDD 5004 5005 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=216970 $D=8
M326 VDD 5012 5013 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=251690 $D=8
M327 VDD 4362 4364 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=252970 $D=8
M328 4758 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=56980 $Y=160970 $D=8
M329 4757 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=56980 $Y=164845 $D=8
M330 5403 4658 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=57195 $Y=112830 $D=8
M331 4346 4348 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=179690 $D=8
M332 4940 4941 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=180970 $D=8
M333 4948 4949 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=215690 $D=8
M334 5004 5005 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=216970 $D=8
M335 5012 5013 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=251690 $D=8
M336 4362 4364 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=252970 $D=8
M337 VDD 4342 4344 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=179690 $D=8
M338 VDD 4938 4939 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=180970 $D=8
M339 VDD 4946 4947 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=215690 $D=8
M340 VDD 5002 5003 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=216970 $D=8
M341 VDD 5010 5011 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=251690 $D=8
M342 VDD 4358 4360 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=252970 $D=8
M343 5402 4657 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=59725 $Y=112830 $D=8
M344 4755 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=60080 $Y=160970 $D=8
M345 4756 948 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=60080 $Y=164845 $D=8
M346 4342 4344 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=179690 $D=8
M347 4938 4939 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=180970 $D=8
M348 4946 4947 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=215690 $D=8
M349 5002 5003 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=216970 $D=8
M350 5010 5011 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=251690 $D=8
M351 4358 4360 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=252970 $D=8
M352 VDD 4546 4548 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=179690 $D=8
M353 VDD 5019 5018 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=180970 $D=8
M354 VDD 5027 5026 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=215690 $D=8
M355 VDD 5083 5082 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=216970 $D=8
M356 VDD 5091 5090 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=251690 $D=8
M357 VDD 5436 5437 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=252970 $D=8
M358 4546 4548 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=179690 $D=8
M359 5019 5018 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=180970 $D=8
M360 5027 5026 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=215690 $D=8
M361 5083 5082 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=216970 $D=8
M362 5091 5090 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=251690 $D=8
M363 5436 5437 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=252970 $D=8
M364 4713 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=67620 $Y=160970 $D=8
M365 4714 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=67620 $Y=164845 $D=8
M366 4869 4664 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=67835 $Y=112830 $D=8
M367 VDD 4542 4544 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=179690 $D=8
M368 VDD 5021 5020 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=180970 $D=8
M369 VDD 5029 5028 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=215690 $D=8
M370 VDD 5085 5084 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=216970 $D=8
M371 VDD 5093 5092 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=251690 $D=8
M372 VDD 5434 5435 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=252970 $D=8
M373 4542 4544 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=179690 $D=8
M374 5021 5020 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=180970 $D=8
M375 5029 5028 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=215690 $D=8
M376 5085 5084 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=216970 $D=8
M377 5093 5092 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=251690 $D=8
M378 5434 5435 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=252970 $D=8
M379 4870 4663 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=70365 $Y=112830 $D=8
M380 4716 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=70720 $Y=160970 $D=8
M381 4715 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=70720 $Y=164845 $D=8
M382 VDD 4538 4540 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=179690 $D=8
M383 VDD 5023 5022 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=180970 $D=8
M384 VDD 5031 5030 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=215690 $D=8
M385 VDD 5087 5086 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=216970 $D=8
M386 VDD 5095 5094 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=251690 $D=8
M387 VDD 5432 5433 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=252970 $D=8
M388 4538 4540 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=179690 $D=8
M389 5023 5022 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=180970 $D=8
M390 5031 5030 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=215690 $D=8
M391 5087 5086 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=216970 $D=8
M392 5095 5094 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=251690 $D=8
M393 5432 5433 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=252970 $D=8
M394 4717 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=73815 $Y=160970 $D=8
M395 4718 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=73815 $Y=164845 $D=8
M396 4871 4662 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=74030 $Y=112830 $D=8
M397 VDD 4534 4536 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=179690 $D=8
M398 VDD 5025 5024 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=180970 $D=8
M399 VDD 5033 5032 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=215690 $D=8
M400 VDD 5089 5088 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=216970 $D=8
M401 VDD 5097 5096 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=251690 $D=8
M402 VDD 5430 5431 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=252970 $D=8
M403 4534 4536 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=179690 $D=8
M404 5025 5024 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=180970 $D=8
M405 5033 5032 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=215690 $D=8
M406 5089 5088 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=216970 $D=8
M407 5097 5096 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=251690 $D=8
M408 5430 5431 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=252970 $D=8
M409 4872 4661 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=76560 $Y=112830 $D=8
M410 4720 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=76915 $Y=160970 $D=8
M411 4719 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=76915 $Y=164845 $D=8
M412 VDD 4282 4284 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=179690 $D=8
M413 VDD 5035 5034 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=180970 $D=8
M414 VDD 5043 5042 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=215690 $D=8
M415 VDD 5099 5098 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=216970 $D=8
M416 VDD 5107 5106 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=251690 $D=8
M417 VDD 5444 5445 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=252970 $D=8
M418 4282 4284 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=179690 $D=8
M419 5035 5034 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=180970 $D=8
M420 5043 5042 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=215690 $D=8
M421 5099 5098 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=216970 $D=8
M422 5107 5106 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=251690 $D=8
M423 5444 5445 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=252970 $D=8
M424 4721 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=80005 $Y=160970 $D=8
M425 4722 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=80005 $Y=164845 $D=8
M426 4873 4660 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=80220 $Y=112830 $D=8
M427 VDD 4278 4280 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=179690 $D=8
M428 VDD 5037 5036 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=180970 $D=8
M429 VDD 5045 5044 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=215690 $D=8
M430 VDD 5101 5100 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=216970 $D=8
M431 VDD 5109 5108 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=251690 $D=8
M432 VDD 5442 5443 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=252970 $D=8
M433 4278 4280 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=179690 $D=8
M434 5037 5036 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=180970 $D=8
M435 5045 5044 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=215690 $D=8
M436 5101 5100 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=216970 $D=8
M437 5109 5108 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=251690 $D=8
M438 5442 5443 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=252970 $D=8
M439 4874 4659 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=82750 $Y=112830 $D=8
M440 4724 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=83105 $Y=160970 $D=8
M441 4723 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=83105 $Y=164845 $D=8
M442 VDD 4290 4292 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=179690 $D=8
M443 VDD 5039 5038 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=180970 $D=8
M444 VDD 5047 5046 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=215690 $D=8
M445 VDD 5103 5102 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=216970 $D=8
M446 VDD 5111 5110 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=251690 $D=8
M447 VDD 5440 5441 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=252970 $D=8
M448 4290 4292 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=179690 $D=8
M449 5039 5038 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=180970 $D=8
M450 5047 5046 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=215690 $D=8
M451 5103 5102 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=216970 $D=8
M452 5111 5110 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=251690 $D=8
M453 5440 5441 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=252970 $D=8
M454 4725 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=86200 $Y=160970 $D=8
M455 4726 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=86200 $Y=164845 $D=8
M456 4875 4658 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=86415 $Y=112830 $D=8
M457 VDD 4286 4288 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=179690 $D=8
M458 VDD 5041 5040 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=180970 $D=8
M459 VDD 5049 5048 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=215690 $D=8
M460 VDD 5105 5104 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=216970 $D=8
M461 VDD 5113 5112 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=251690 $D=8
M462 VDD 5438 5439 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=252970 $D=8
M463 4286 4288 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=179690 $D=8
M464 5041 5040 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=180970 $D=8
M465 5049 5048 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=215690 $D=8
M466 5105 5104 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=216970 $D=8
M467 5113 5112 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=251690 $D=8
M468 5438 5439 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=252970 $D=8
M469 4819 4657 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=88945 $Y=112830 $D=8
M470 940 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=89120 $Y=160970 $D=8
M471 941 4219 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=89120 $Y=164845 $D=8
M472 953 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=92575 $Y=160970 $D=8
M473 954 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=92575 $Y=164845 $D=8
M474 VDD 4562 4564 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=179690 $D=8
M475 VDD 5056 5057 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=180970 $D=8
M476 VDD 5064 5065 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=215690 $D=8
M477 VDD 5120 5121 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=216970 $D=8
M478 VDD 5128 5129 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=251690 $D=8
M479 VDD 5452 5453 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=252970 $D=8
M480 4823 4664 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=92620 $Y=112830 $D=8
M481 4562 4564 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=179690 $D=8
M482 5056 5057 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=180970 $D=8
M483 5064 5065 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=215690 $D=8
M484 5120 5121 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=216970 $D=8
M485 5128 5129 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=251690 $D=8
M486 5452 5453 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=252970 $D=8
M487 5415 4663 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=95145 $Y=112830 $D=8
M488 4797 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=95500 $Y=160970 $D=8
M489 4798 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=95500 $Y=164845 $D=8
M490 VDD 4558 4560 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=179690 $D=8
M491 VDD 5054 5055 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=180970 $D=8
M492 VDD 5062 5063 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=215690 $D=8
M493 VDD 5118 5119 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=216970 $D=8
M494 VDD 5126 5127 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=251690 $D=8
M495 VDD 5450 5451 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=252970 $D=8
M496 4558 4560 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=179690 $D=8
M497 5054 5055 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=180970 $D=8
M498 5062 5063 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=215690 $D=8
M499 5118 5119 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=216970 $D=8
M500 5126 5127 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=251690 $D=8
M501 5450 5451 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=252970 $D=8
M502 4796 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=98595 $Y=160970 $D=8
M503 4795 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=98595 $Y=164845 $D=8
M504 VDD 4554 4556 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=179690 $D=8
M505 VDD 5052 5053 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=180970 $D=8
M506 VDD 5060 5061 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=215690 $D=8
M507 VDD 5116 5117 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=216970 $D=8
M508 VDD 5124 5125 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=251690 $D=8
M509 VDD 5448 5449 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=252970 $D=8
M510 5414 4662 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=98810 $Y=112830 $D=8
M511 4554 4556 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=179690 $D=8
M512 5052 5053 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=180970 $D=8
M513 5060 5061 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=215690 $D=8
M514 5116 5117 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=216970 $D=8
M515 5124 5125 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=251690 $D=8
M516 5448 5449 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=252970 $D=8
M517 5413 4661 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=101340 $Y=112830 $D=8
M518 4793 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=101695 $Y=160970 $D=8
M519 4794 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=101695 $Y=164845 $D=8
M520 VDD 4550 4552 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=179690 $D=8
M521 VDD 5050 5051 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=180970 $D=8
M522 VDD 5058 5059 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=215690 $D=8
M523 VDD 5114 5115 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=216970 $D=8
M524 VDD 5122 5123 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=251690 $D=8
M525 VDD 5446 5447 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=252970 $D=8
M526 4550 4552 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=179690 $D=8
M527 5050 5051 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=180970 $D=8
M528 5058 5059 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=215690 $D=8
M529 5114 5115 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=216970 $D=8
M530 5122 5123 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=251690 $D=8
M531 5446 5447 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=252970 $D=8
M532 VDD 4386 4388 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=179690 $D=8
M533 VDD 5072 5073 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=180970 $D=8
M534 VDD 5080 5081 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=215690 $D=8
M535 VDD 5136 5137 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=216970 $D=8
M536 VDD 5144 5145 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=251690 $D=8
M537 VDD 5460 5461 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=252970 $D=8
M538 4770 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=104785 $Y=160970 $D=8
M539 4769 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=104785 $Y=164845 $D=8
M540 5412 4660 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=105000 $Y=112830 $D=8
M541 4386 4388 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=179690 $D=8
M542 5072 5073 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=180970 $D=8
M543 5080 5081 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=215690 $D=8
M544 5136 5137 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=216970 $D=8
M545 5144 5145 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=251690 $D=8
M546 5460 5461 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=252970 $D=8
M547 5411 4659 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=107530 $Y=112830 $D=8
M548 VDD 4382 4384 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=179690 $D=8
M549 VDD 5070 5071 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=180970 $D=8
M550 VDD 5078 5079 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=215690 $D=8
M551 VDD 5134 5135 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=216970 $D=8
M552 VDD 5142 5143 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=251690 $D=8
M553 VDD 5458 5459 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=252970 $D=8
M554 4767 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=107885 $Y=160970 $D=8
M555 4768 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=107885 $Y=164845 $D=8
M556 4382 4384 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=179690 $D=8
M557 5070 5071 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=180970 $D=8
M558 5078 5079 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=215690 $D=8
M559 5134 5135 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=216970 $D=8
M560 5142 5143 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=251690 $D=8
M561 5458 5459 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=252970 $D=8
M562 VDD 4378 4380 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=179690 $D=8
M563 VDD 5068 5069 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=180970 $D=8
M564 VDD 5076 5077 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=215690 $D=8
M565 VDD 5132 5133 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=216970 $D=8
M566 VDD 5140 5141 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=251690 $D=8
M567 VDD 5456 5457 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=252970 $D=8
M568 4766 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=110980 $Y=160970 $D=8
M569 4765 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=110980 $Y=164845 $D=8
M570 5410 4658 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=111195 $Y=112830 $D=8
M571 4378 4380 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=179690 $D=8
M572 5068 5069 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=180970 $D=8
M573 5076 5077 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=215690 $D=8
M574 5132 5133 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=216970 $D=8
M575 5140 5141 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=251690 $D=8
M576 5456 5457 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=252970 $D=8
M577 VDD 4374 4376 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=179690 $D=8
M578 VDD 5066 5067 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=180970 $D=8
M579 VDD 5074 5075 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=215690 $D=8
M580 VDD 5130 5131 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=216970 $D=8
M581 VDD 5138 5139 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=251690 $D=8
M582 VDD 5454 5455 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=252970 $D=8
M583 5409 4657 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=113725 $Y=112830 $D=8
M584 4763 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=114080 $Y=160970 $D=8
M585 4764 952 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=114080 $Y=164845 $D=8
M586 4374 4376 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=179690 $D=8
M587 5066 5067 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=180970 $D=8
M588 5074 5075 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=215690 $D=8
M589 5130 5131 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=216970 $D=8
M590 5138 5139 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=251690 $D=8
M591 5454 5455 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=252970 $D=8
M592 VDD 4645 4646 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=179690 $D=8
M593 VDD 5494 5495 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=180970 $D=8
M594 VDD 5496 5497 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=188690 $D=8
M595 VDD 5498 5499 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=189970 $D=8
M596 VDD 5500 5501 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=197690 $D=8
M597 VDD 5502 5503 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=198970 $D=8
M598 VDD 5504 5505 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=206690 $D=8
M599 VDD 5506 5507 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=207970 $D=8
M600 VDD 5508 5509 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=215690 $D=8
M601 VDD 5510 5511 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=216970 $D=8
M602 VDD 5512 5513 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=224690 $D=8
M603 VDD 5514 5515 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=225970 $D=8
M604 VDD 5516 5517 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=233690 $D=8
M605 VDD 5518 5519 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=234970 $D=8
M606 VDD 5520 5521 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=242690 $D=8
M607 VDD 5522 5523 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=243970 $D=8
M608 VDD 5524 5525 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=251690 $D=8
M609 VDD 4647 4648 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=252970 $D=8
M610 VDD VSS VDD VDD pfet_05v0 L=2.365e-06 W=8.19e-05 AD=0 AS=6.1309e-11 PD=0 PS=0.000217698 NRD=0 NRS=11.8457 m=1 nf=36 $X=10835 $Y=171065 $D=8
M611 4645 4646 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=179690 $D=8
M612 5494 5495 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=180970 $D=8
M613 5496 5497 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=188690 $D=8
M614 5498 5499 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=189970 $D=8
M615 5500 5501 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=197690 $D=8
M616 5502 5503 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=198970 $D=8
M617 5504 5505 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=206690 $D=8
M618 5506 5507 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=207970 $D=8
M619 5508 5509 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=215690 $D=8
M620 5510 5511 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=216970 $D=8
M621 5512 5513 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=224690 $D=8
M622 5514 5515 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=225970 $D=8
M623 5516 5517 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=233690 $D=8
M624 5518 5519 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=234970 $D=8
M625 5520 5521 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=242690 $D=8
M626 5522 5523 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=243970 $D=8
M627 5524 5525 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=251690 $D=8
M628 4647 4648 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=252970 $D=8
M629 VDD VSS VDD VDD pfet_05v0 L=3.94e-06 W=9.3415e-05 AD=0 AS=5.61039e-11 PD=0 PS=0.00021824 NRD=0 NRS=1.85805 m=1 nf=17 $X=146370 $Y=180915 $D=8
M630 VDD 4854 4222 VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=156680 $Y=180895 $D=8
M631 4229 4856 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=213535 $D=8
M632 VDD 4858 4230 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=216895 $D=8
M633 4237 4860 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=156680 $Y=249535 $D=8
M634 4827 VDD VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=180895 $D=8
M635 VDD 918 4827 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=182015 $D=8
M636 4827 926 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=183135 $D=8
M637 VDD 919 4829 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=213535 $D=8
M638 4829 918 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=214655 $D=8
M639 VDD VDD 4829 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=215775 $D=8
M640 4831 VDD VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=216895 $D=8
M641 VDD 917 4831 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=218015 $D=8
M642 4831 926 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=219135 $D=8
M643 VDD 919 4833 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=249535 $D=8
M644 4833 917 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=250655 $D=8
M645 VDD VDD 4833 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=251775 $D=8
M646 4817 1 VDD VDD pfet_05v0 L=5.95e-07 W=2.28e-06 AD=5.985e-13 AS=1.3566e-12 PD=2.805e-06 PS=5.75e-06 NRD=0.115132 NRS=0.260965 m=1 nf=1 $X=233770 $Y=57780 $D=8
M647 617 787 VDD VDD pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=233770 $Y=63100 $D=8
M648 787 CLK 4817 VDD pfet_05v0 L=5.95e-07 W=2.28e-06 AD=1.3566e-12 AS=5.985e-13 PD=5.75e-06 PS=2.805e-06 NRD=0.260965 NRS=0.115132 m=1 nf=1 $X=234890 $Y=57780 $D=8
M649 616 619 VDD VDD pfet_05v0 L=6e-07 W=1.134e-05 AD=2.9484e-12 AS=4.9896e-12 PD=1.238e-05 PS=2.444e-05 NRD=0.0917108 NRS=0.155203 m=1 nf=2 $X=242235 $Y=57810 $D=8
M650 281 865 VDD VDD pfet_05v0 L=1e-06 W=9e-07 AD=3.96e-13 AS=3.96e-13 PD=2.68e-06 PS=2.68e-06 NRD=0.488889 NRS=0.488889 m=1 nf=1 $X=243265 $Y=42525 $D=8
M651 CEN 617 619 VDD pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=245925 $Y=59010 $D=8
M652 618 787 619 VDD pfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=245925 $Y=64875 $D=8
M653 317 281 VDD VDD pfet_05v0 L=6e-07 W=1.89e-06 AD=8.316e-13 AS=8.316e-13 PD=4.66e-06 PS=4.66e-06 NRD=0.232804 NRS=0.232804 m=1 nf=1 $X=246495 $Y=41535 $D=8
M654 354 317 VDD VDD pfet_05v0 L=6e-07 W=7.54e-06 AD=1.9604e-12 AS=3.3176e-12 PD=8.58e-06 PS=1.684e-05 NRD=0.137931 NRS=0.233422 m=1 nf=2 $X=249065 $Y=39655 $D=8
M655 250 468 VDD VDD pfet_05v0 L=6e-07 W=0.0001248 AD=3.2448e-11 AS=3.69283e-11 PD=0.00013 PS=0.000130718 NRD=0.208333 NRS=0.237099 m=1 nf=10 $X=240535 $Y=94430 $D=8
M656 445 354 VDD VDD pfet_05v0 L=6e-07 W=1.95e-05 AD=5.07e-12 AS=8.58e-12 PD=2.002e-05 PS=3.988e-05 NRD=0.0133333 NRS=0.0225641 m=1 nf=1 $X=256125 $Y=53590 $D=8
M657 VDD CLK 445 VDD pfet_05v0 L=6e-07 W=1.95e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=257245 $Y=53590 $D=8
M658 445 616 VDD VDD pfet_05v0 L=6e-07 W=1.95e-05 AD=8.58e-12 AS=5.07e-12 PD=3.988e-05 PS=2.002e-05 NRD=0.0225641 NRS=0.0133333 m=1 nf=1 $X=258365 $Y=53590 $D=8
M659 VDD 495 468 VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=9.9792e-12 PD=2.32e-05 PS=4.624e-05 NRD=0.0114638 NRS=0.0194004 m=1 nf=1 $X=262120 $Y=50420 $D=8
M660 468 445 VDD VDD pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.64e-05 PS=4.64e-05 NRD=0.0229277 NRS=0.0229277 m=1 nf=2 $X=263240 $Y=50420 $D=8
M661 468 495 VDD VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=9.9792e-12 AS=5.8968e-12 PD=4.624e-05 PS=2.32e-05 NRD=0.0194004 NRS=0.0114638 m=1 nf=1 $X=265480 $Y=50420 $D=8
M662 VDD 4855 4238 VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=258945 $Y=180895 $D=8
M663 4245 4857 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=213535 $D=8
M664 VDD 4859 4246 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=216895 $D=8
M665 4253 4861 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=258945 $Y=249535 $D=8
M666 VDD 468 495 VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=9.9792e-12 PD=2.32e-05 PS=4.624e-05 NRD=0.0114638 NRS=0.0194004 m=1 nf=1 $X=268545 $Y=50420 $D=8
M667 495 607 VDD VDD pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.64e-05 PS=4.64e-05 NRD=0.0229277 NRS=0.0229277 m=1 nf=2 $X=269665 $Y=50420 $D=8
M668 495 468 VDD VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=9.9792e-12 AS=5.8968e-12 PD=4.624e-05 PS=2.32e-05 NRD=0.0194004 NRS=0.0114638 m=1 nf=1 $X=271905 $Y=50420 $D=8
M669 1 250 VDD VDD pfet_05v0 L=6e-07 W=0.0003674 AD=9.5524e-11 AS=1.02119e-10 PD=0.0003778 PS=0.000378518 NRD=0.28307 NRS=0.302613 m=1 nf=20 $X=253180 $Y=88540 $D=8
M670 VDD VSS VDD VDD pfet_05v0 L=3.94e-06 W=9.3415e-05 AD=0 AS=5.61039e-11 PD=0 PS=0.00021824 NRD=0 NRS=1.85805 m=1 nf=17 $X=273750 $Y=180915 $D=8
M671 VDD 4649 4650 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=179690 $D=8
M672 VDD 5534 5536 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=180970 $D=8
M673 VDD 5535 5537 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=188690 $D=8
M674 VDD 5538 5540 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=189970 $D=8
M675 VDD 5539 5541 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=197690 $D=8
M676 VDD 5542 5544 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=198970 $D=8
M677 VDD 5543 5545 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=206690 $D=8
M678 VDD 5546 5548 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=207970 $D=8
M679 VDD 5547 5549 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=215690 $D=8
M680 VDD 5550 5552 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=216970 $D=8
M681 VDD 5551 5553 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=224690 $D=8
M682 VDD 5554 5556 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=225970 $D=8
M683 VDD 5555 5557 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=233690 $D=8
M684 VDD 5558 5560 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=234970 $D=8
M685 VDD 5559 5561 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=242690 $D=8
M686 VDD 5562 5564 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=243970 $D=8
M687 VDD 5563 5565 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=251690 $D=8
M688 VDD 4651 4652 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=252970 $D=8
M689 4649 4650 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=179690 $D=8
M690 5534 5536 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=180970 $D=8
M691 5535 5537 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=188690 $D=8
M692 5538 5540 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=189970 $D=8
M693 5539 5541 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=197690 $D=8
M694 5542 5544 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=198970 $D=8
M695 5543 5545 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=206690 $D=8
M696 5546 5548 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=207970 $D=8
M697 5547 5549 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=215690 $D=8
M698 5550 5552 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=216970 $D=8
M699 5551 5553 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=224690 $D=8
M700 5554 5556 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=225970 $D=8
M701 5555 5557 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=233690 $D=8
M702 5558 5560 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=234970 $D=8
M703 5559 5561 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=242690 $D=8
M704 5562 5564 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=243970 $D=8
M705 5563 5565 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=251690 $D=8
M706 4651 4652 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=252970 $D=8
M707 VDD 4578 4580 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=179690 $D=8
M708 VDD 5147 5146 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=180970 $D=8
M709 VDD 5155 5154 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=215690 $D=8
M710 VDD 5211 5210 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=216970 $D=8
M711 VDD 5219 5218 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=251690 $D=8
M712 VDD 4402 4404 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=252970 $D=8
M713 4578 4580 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=179690 $D=8
M714 5147 5146 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=180970 $D=8
M715 5155 5154 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=215690 $D=8
M716 5211 5210 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=216970 $D=8
M717 5219 5218 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=251690 $D=8
M718 4402 4404 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=252970 $D=8
M719 4727 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=311500 $Y=160970 $D=8
M720 4728 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=311500 $Y=164845 $D=8
M721 4876 4666 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=311715 $Y=112830 $D=8
M722 VDD 4574 4576 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=179690 $D=8
M723 VDD 5149 5148 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=180970 $D=8
M724 VDD 5157 5156 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=215690 $D=8
M725 VDD 5213 5212 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=216970 $D=8
M726 VDD 5221 5220 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=251690 $D=8
M727 VDD 4398 4400 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=252970 $D=8
M728 4574 4576 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=179690 $D=8
M729 5149 5148 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=180970 $D=8
M730 5157 5156 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=215690 $D=8
M731 5213 5212 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=216970 $D=8
M732 5221 5220 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=251690 $D=8
M733 4398 4400 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=252970 $D=8
M734 4877 4667 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=314245 $Y=112830 $D=8
M735 4730 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=314600 $Y=160970 $D=8
M736 4729 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=314600 $Y=164845 $D=8
M737 VDD 4570 4572 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=179690 $D=8
M738 VDD 5151 5150 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=180970 $D=8
M739 VDD 5159 5158 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=215690 $D=8
M740 VDD 5215 5214 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=216970 $D=8
M741 VDD 5223 5222 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=251690 $D=8
M742 VDD 4394 4396 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=252970 $D=8
M743 4570 4572 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=179690 $D=8
M744 5151 5150 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=180970 $D=8
M745 5159 5158 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=215690 $D=8
M746 5215 5214 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=216970 $D=8
M747 5223 5222 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=251690 $D=8
M748 4394 4396 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=252970 $D=8
M749 4731 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=317695 $Y=160970 $D=8
M750 4732 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=317695 $Y=164845 $D=8
M751 4878 4668 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=317910 $Y=112830 $D=8
M752 VDD 4566 4568 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=179690 $D=8
M753 VDD 5153 5152 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=180970 $D=8
M754 VDD 5161 5160 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=215690 $D=8
M755 VDD 5217 5216 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=216970 $D=8
M756 VDD 5225 5224 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=251690 $D=8
M757 VDD 4390 4392 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=252970 $D=8
M758 4566 4568 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=179690 $D=8
M759 5153 5152 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=180970 $D=8
M760 5161 5160 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=215690 $D=8
M761 5217 5216 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=216970 $D=8
M762 5225 5224 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=251690 $D=8
M763 4390 4392 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=252970 $D=8
M764 4879 4669 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=320440 $Y=112830 $D=8
M765 4734 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=320795 $Y=160970 $D=8
M766 4733 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=320795 $Y=164845 $D=8
M767 VDD 4298 4300 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=179690 $D=8
M768 VDD 5163 5162 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=180970 $D=8
M769 VDD 5171 5170 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=215690 $D=8
M770 VDD 5227 5226 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=216970 $D=8
M771 VDD 5235 5234 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=251690 $D=8
M772 VDD 4418 4420 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=252970 $D=8
M773 4298 4300 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=179690 $D=8
M774 5163 5162 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=180970 $D=8
M775 5171 5170 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=215690 $D=8
M776 5227 5226 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=216970 $D=8
M777 5235 5234 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=251690 $D=8
M778 4418 4420 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=252970 $D=8
M779 4735 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=323885 $Y=160970 $D=8
M780 4736 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=323885 $Y=164845 $D=8
M781 4880 4670 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=324100 $Y=112830 $D=8
M782 VDD 4294 4296 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=179690 $D=8
M783 VDD 5165 5164 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=180970 $D=8
M784 VDD 5173 5172 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=215690 $D=8
M785 VDD 5229 5228 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=216970 $D=8
M786 VDD 5237 5236 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=251690 $D=8
M787 VDD 4414 4416 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=252970 $D=8
M788 4294 4296 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=179690 $D=8
M789 5165 5164 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=180970 $D=8
M790 5173 5172 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=215690 $D=8
M791 5229 5228 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=216970 $D=8
M792 5237 5236 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=251690 $D=8
M793 4414 4416 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=252970 $D=8
M794 4881 4671 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=326630 $Y=112830 $D=8
M795 4738 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=326985 $Y=160970 $D=8
M796 4737 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=326985 $Y=164845 $D=8
M797 VDD 4306 4308 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=179690 $D=8
M798 VDD 5167 5166 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=180970 $D=8
M799 VDD 5175 5174 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=215690 $D=8
M800 VDD 5231 5230 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=216970 $D=8
M801 VDD 5239 5238 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=251690 $D=8
M802 VDD 4410 4412 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=252970 $D=8
M803 4306 4308 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=179690 $D=8
M804 5167 5166 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=180970 $D=8
M805 5175 5174 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=215690 $D=8
M806 5231 5230 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=216970 $D=8
M807 5239 5238 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=251690 $D=8
M808 4410 4412 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=252970 $D=8
M809 4739 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=330080 $Y=160970 $D=8
M810 4740 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=330080 $Y=164845 $D=8
M811 4882 4672 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=330295 $Y=112830 $D=8
M812 VDD 4302 4304 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=179690 $D=8
M813 VDD 5169 5168 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=180970 $D=8
M814 VDD 5177 5176 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=215690 $D=8
M815 VDD 5233 5232 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=216970 $D=8
M816 VDD 5241 5240 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=251690 $D=8
M817 VDD 4406 4408 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=252970 $D=8
M818 4302 4304 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=179690 $D=8
M819 5169 5168 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=180970 $D=8
M820 5177 5176 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=215690 $D=8
M821 5233 5232 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=216970 $D=8
M822 5241 5240 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=251690 $D=8
M823 4406 4408 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=252970 $D=8
M824 4820 4673 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=332825 $Y=112830 $D=8
M825 943 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=333000 $Y=160970 $D=8
M826 944 4220 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=333000 $Y=164845 $D=8
M827 957 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=336455 $Y=160970 $D=8
M828 958 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=336455 $Y=164845 $D=8
M829 VDD 4594 4596 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=179690 $D=8
M830 VDD 5184 5185 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=180970 $D=8
M831 VDD 5192 5193 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=215690 $D=8
M832 VDD 5248 5249 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=216970 $D=8
M833 VDD 5256 5257 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=251690 $D=8
M834 VDD 4610 4612 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=252970 $D=8
M835 4824 4666 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=336500 $Y=112830 $D=8
M836 4594 4596 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=179690 $D=8
M837 5184 5185 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=180970 $D=8
M838 5192 5193 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=215690 $D=8
M839 5248 5249 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=216970 $D=8
M840 5256 5257 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=251690 $D=8
M841 4610 4612 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=252970 $D=8
M842 5422 4667 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=339025 $Y=112830 $D=8
M843 4803 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=339380 $Y=160970 $D=8
M844 4804 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=339380 $Y=164845 $D=8
M845 VDD 4590 4592 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=179690 $D=8
M846 VDD 5182 5183 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=180970 $D=8
M847 VDD 5190 5191 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=215690 $D=8
M848 VDD 5246 5247 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=216970 $D=8
M849 VDD 5254 5255 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=251690 $D=8
M850 VDD 4606 4608 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=252970 $D=8
M851 4590 4592 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=179690 $D=8
M852 5182 5183 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=180970 $D=8
M853 5190 5191 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=215690 $D=8
M854 5246 5247 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=216970 $D=8
M855 5254 5255 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=251690 $D=8
M856 4606 4608 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=252970 $D=8
M857 4802 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=342475 $Y=160970 $D=8
M858 4801 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=342475 $Y=164845 $D=8
M859 VDD 4586 4588 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=179690 $D=8
M860 VDD 5180 5181 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=180970 $D=8
M861 VDD 5188 5189 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=215690 $D=8
M862 VDD 5244 5245 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=216970 $D=8
M863 VDD 5252 5253 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=251690 $D=8
M864 VDD 4602 4604 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=252970 $D=8
M865 5421 4668 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=342690 $Y=112830 $D=8
M866 4586 4588 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=179690 $D=8
M867 5180 5181 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=180970 $D=8
M868 5188 5189 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=215690 $D=8
M869 5244 5245 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=216970 $D=8
M870 5252 5253 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=251690 $D=8
M871 4602 4604 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=252970 $D=8
M872 5420 4669 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=345220 $Y=112830 $D=8
M873 4799 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=345575 $Y=160970 $D=8
M874 4800 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=345575 $Y=164845 $D=8
M875 VDD 4582 4584 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=179690 $D=8
M876 VDD 5178 5179 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=180970 $D=8
M877 VDD 5186 5187 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=215690 $D=8
M878 VDD 5242 5243 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=216970 $D=8
M879 VDD 5250 5251 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=251690 $D=8
M880 VDD 4598 4600 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=252970 $D=8
M881 4582 4584 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=179690 $D=8
M882 5178 5179 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=180970 $D=8
M883 5186 5187 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=215690 $D=8
M884 5242 5243 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=216970 $D=8
M885 5250 5251 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=251690 $D=8
M886 4598 4600 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=252970 $D=8
M887 VDD 4434 4436 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=179690 $D=8
M888 VDD 5200 5201 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=180970 $D=8
M889 VDD 5208 5209 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=215690 $D=8
M890 VDD 5264 5265 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=216970 $D=8
M891 VDD 5272 5273 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=251690 $D=8
M892 VDD 4450 4452 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=252970 $D=8
M893 4778 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=348665 $Y=160970 $D=8
M894 4777 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=348665 $Y=164845 $D=8
M895 5419 4670 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=348880 $Y=112830 $D=8
M896 4434 4436 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=179690 $D=8
M897 5200 5201 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=180970 $D=8
M898 5208 5209 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=215690 $D=8
M899 5264 5265 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=216970 $D=8
M900 5272 5273 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=251690 $D=8
M901 4450 4452 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=252970 $D=8
M902 5418 4671 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=351410 $Y=112830 $D=8
M903 VDD 4430 4432 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=179690 $D=8
M904 VDD 5198 5199 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=180970 $D=8
M905 VDD 5206 5207 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=215690 $D=8
M906 VDD 5262 5263 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=216970 $D=8
M907 VDD 5270 5271 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=251690 $D=8
M908 VDD 4446 4448 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=252970 $D=8
M909 4775 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=351765 $Y=160970 $D=8
M910 4776 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=351765 $Y=164845 $D=8
M911 4430 4432 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=179690 $D=8
M912 5198 5199 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=180970 $D=8
M913 5206 5207 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=215690 $D=8
M914 5262 5263 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=216970 $D=8
M915 5270 5271 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=251690 $D=8
M916 4446 4448 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=252970 $D=8
M917 VDD 4426 4428 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=179690 $D=8
M918 VDD 5196 5197 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=180970 $D=8
M919 VDD 5204 5205 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=215690 $D=8
M920 VDD 5260 5261 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=216970 $D=8
M921 VDD 5268 5269 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=251690 $D=8
M922 VDD 4442 4444 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=252970 $D=8
M923 4774 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=354860 $Y=160970 $D=8
M924 4773 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=354860 $Y=164845 $D=8
M925 5417 4672 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=355075 $Y=112830 $D=8
M926 4426 4428 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=179690 $D=8
M927 5196 5197 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=180970 $D=8
M928 5204 5205 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=215690 $D=8
M929 5260 5261 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=216970 $D=8
M930 5268 5269 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=251690 $D=8
M931 4442 4444 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=252970 $D=8
M932 VDD 4422 4424 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=179690 $D=8
M933 VDD 5194 5195 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=180970 $D=8
M934 VDD 5202 5203 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=215690 $D=8
M935 VDD 5258 5259 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=216970 $D=8
M936 VDD 5266 5267 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=251690 $D=8
M937 VDD 4438 4440 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=252970 $D=8
M938 5416 4673 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=357605 $Y=112830 $D=8
M939 4771 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=357960 $Y=160970 $D=8
M940 4772 955 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=357960 $Y=164845 $D=8
M941 4422 4424 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=179690 $D=8
M942 5194 5195 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=180970 $D=8
M943 5202 5203 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=215690 $D=8
M944 5258 5259 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=216970 $D=8
M945 5266 5267 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=251690 $D=8
M946 4438 4440 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=252970 $D=8
M947 VDD 4626 4628 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=179690 $D=8
M948 VDD 5275 5274 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=180970 $D=8
M949 VDD 5283 5282 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=215690 $D=8
M950 VDD 5339 5338 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=216970 $D=8
M951 VDD 5347 5346 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=251690 $D=8
M952 VDD 5468 5469 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=252970 $D=8
M953 4626 4628 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=179690 $D=8
M954 5275 5274 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=180970 $D=8
M955 5283 5282 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=215690 $D=8
M956 5339 5338 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=216970 $D=8
M957 5347 5346 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=251690 $D=8
M958 5468 5469 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=252970 $D=8
M959 4741 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=365500 $Y=160970 $D=8
M960 4742 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=365500 $Y=164845 $D=8
M961 4883 4666 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=365715 $Y=112830 $D=8
M962 VDD 4622 4624 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=179690 $D=8
M963 VDD 5277 5276 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=180970 $D=8
M964 VDD 5285 5284 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=215690 $D=8
M965 VDD 5341 5340 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=216970 $D=8
M966 VDD 5349 5348 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=251690 $D=8
M967 VDD 5466 5467 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=252970 $D=8
M968 4622 4624 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=179690 $D=8
M969 5277 5276 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=180970 $D=8
M970 5285 5284 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=215690 $D=8
M971 5341 5340 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=216970 $D=8
M972 5349 5348 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=251690 $D=8
M973 5466 5467 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=252970 $D=8
M974 4884 4667 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=368245 $Y=112830 $D=8
M975 4744 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=368600 $Y=160970 $D=8
M976 4743 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=368600 $Y=164845 $D=8
M977 VDD 4618 4620 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=179690 $D=8
M978 VDD 5279 5278 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=180970 $D=8
M979 VDD 5287 5286 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=215690 $D=8
M980 VDD 5343 5342 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=216970 $D=8
M981 VDD 5351 5350 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=251690 $D=8
M982 VDD 5464 5465 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=252970 $D=8
M983 4618 4620 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=179690 $D=8
M984 5279 5278 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=180970 $D=8
M985 5287 5286 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=215690 $D=8
M986 5343 5342 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=216970 $D=8
M987 5351 5350 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=251690 $D=8
M988 5464 5465 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=252970 $D=8
M989 4745 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=371695 $Y=160970 $D=8
M990 4746 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=371695 $Y=164845 $D=8
M991 4885 4668 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=371910 $Y=112830 $D=8
M992 VDD 4614 4616 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=179690 $D=8
M993 VDD 5281 5280 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=180970 $D=8
M994 VDD 5289 5288 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=215690 $D=8
M995 VDD 5345 5344 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=216970 $D=8
M996 VDD 5353 5352 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=251690 $D=8
M997 VDD 5462 5463 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=252970 $D=8
M998 4614 4616 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=179690 $D=8
M999 5281 5280 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=180970 $D=8
M1000 5289 5288 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=215690 $D=8
M1001 5345 5344 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=216970 $D=8
M1002 5353 5352 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=251690 $D=8
M1003 5462 5463 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=252970 $D=8
M1004 4886 4669 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=374440 $Y=112830 $D=8
M1005 4748 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=374795 $Y=160970 $D=8
M1006 4747 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=374795 $Y=164845 $D=8
M1007 VDD 4314 4316 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=179690 $D=8
M1008 VDD 5291 5290 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=180970 $D=8
M1009 VDD 5299 5298 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=215690 $D=8
M1010 VDD 5355 5354 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=216970 $D=8
M1011 VDD 5363 5362 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=251690 $D=8
M1012 VDD 5476 5477 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=252970 $D=8
M1013 4314 4316 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=179690 $D=8
M1014 5291 5290 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=180970 $D=8
M1015 5299 5298 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=215690 $D=8
M1016 5355 5354 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=216970 $D=8
M1017 5363 5362 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=251690 $D=8
M1018 5476 5477 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=252970 $D=8
M1019 4749 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=377885 $Y=160970 $D=8
M1020 4750 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=377885 $Y=164845 $D=8
M1021 4887 4670 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=378100 $Y=112830 $D=8
M1022 VDD 4310 4312 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=179690 $D=8
M1023 VDD 5293 5292 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=180970 $D=8
M1024 VDD 5301 5300 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=215690 $D=8
M1025 VDD 5357 5356 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=216970 $D=8
M1026 VDD 5365 5364 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=251690 $D=8
M1027 VDD 5474 5475 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=252970 $D=8
M1028 4310 4312 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=179690 $D=8
M1029 5293 5292 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=180970 $D=8
M1030 5301 5300 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=215690 $D=8
M1031 5357 5356 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=216970 $D=8
M1032 5365 5364 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=251690 $D=8
M1033 5474 5475 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=252970 $D=8
M1034 4888 4671 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=380630 $Y=112830 $D=8
M1035 4752 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=380985 $Y=160970 $D=8
M1036 4751 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=380985 $Y=164845 $D=8
M1037 VDD 4322 4324 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=179690 $D=8
M1038 VDD 5295 5294 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=180970 $D=8
M1039 VDD 5303 5302 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=215690 $D=8
M1040 VDD 5359 5358 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=216970 $D=8
M1041 VDD 5367 5366 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=251690 $D=8
M1042 VDD 5472 5473 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=252970 $D=8
M1043 4322 4324 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=179690 $D=8
M1044 5295 5294 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=180970 $D=8
M1045 5303 5302 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=215690 $D=8
M1046 5359 5358 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=216970 $D=8
M1047 5367 5366 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=251690 $D=8
M1048 5472 5473 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=252970 $D=8
M1049 4753 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=384080 $Y=160970 $D=8
M1050 4754 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=384080 $Y=164845 $D=8
M1051 4889 4672 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=384295 $Y=112830 $D=8
M1052 VDD 4318 4320 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=179690 $D=8
M1053 VDD 5297 5296 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=180970 $D=8
M1054 VDD 5305 5304 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=215690 $D=8
M1055 VDD 5361 5360 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=216970 $D=8
M1056 VDD 5369 5368 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=251690 $D=8
M1057 VDD 5470 5471 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=252970 $D=8
M1058 4318 4320 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=179690 $D=8
M1059 5297 5296 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=180970 $D=8
M1060 5305 5304 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=215690 $D=8
M1061 5361 5360 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=216970 $D=8
M1062 5369 5368 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=251690 $D=8
M1063 5470 5471 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=252970 $D=8
M1064 4821 4673 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=386825 $Y=112830 $D=8
M1065 946 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=387000 $Y=160970 $D=8
M1066 947 4221 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=387000 $Y=164845 $D=8
M1067 960 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=390455 $Y=160970 $D=8
M1068 961 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=390455 $Y=164845 $D=8
M1069 VDD 4642 4644 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=179690 $D=8
M1070 VDD 5312 5313 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=180970 $D=8
M1071 VDD 5320 5321 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=215690 $D=8
M1072 VDD 5376 5377 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=216970 $D=8
M1073 VDD 5384 5385 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=251690 $D=8
M1074 VDD 5484 5485 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=252970 $D=8
M1075 4825 4666 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=390500 $Y=112830 $D=8
M1076 4642 4644 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=179690 $D=8
M1077 5312 5313 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=180970 $D=8
M1078 5320 5321 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=215690 $D=8
M1079 5376 5377 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=216970 $D=8
M1080 5384 5385 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=251690 $D=8
M1081 5484 5485 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=252970 $D=8
M1082 5429 4667 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=393025 $Y=112830 $D=8
M1083 4809 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=393380 $Y=160970 $D=8
M1084 4810 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=393380 $Y=164845 $D=8
M1085 VDD 4638 4640 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=179690 $D=8
M1086 VDD 5310 5311 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=180970 $D=8
M1087 VDD 5318 5319 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=215690 $D=8
M1088 VDD 5374 5375 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=216970 $D=8
M1089 VDD 5382 5383 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=251690 $D=8
M1090 VDD 5482 5483 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=252970 $D=8
M1091 4638 4640 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=179690 $D=8
M1092 5310 5311 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=180970 $D=8
M1093 5318 5319 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=215690 $D=8
M1094 5374 5375 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=216970 $D=8
M1095 5382 5383 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=251690 $D=8
M1096 5482 5483 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=252970 $D=8
M1097 4808 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=396475 $Y=160970 $D=8
M1098 4807 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=396475 $Y=164845 $D=8
M1099 VDD 4634 4636 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=179690 $D=8
M1100 VDD 5308 5309 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=180970 $D=8
M1101 VDD 5316 5317 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=215690 $D=8
M1102 VDD 5372 5373 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=216970 $D=8
M1103 VDD 5380 5381 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=251690 $D=8
M1104 VDD 5480 5481 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=252970 $D=8
M1105 5428 4668 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=396690 $Y=112830 $D=8
M1106 4634 4636 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=179690 $D=8
M1107 5308 5309 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=180970 $D=8
M1108 5316 5317 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=215690 $D=8
M1109 5372 5373 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=216970 $D=8
M1110 5380 5381 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=251690 $D=8
M1111 5480 5481 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=252970 $D=8
M1112 5427 4669 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=399220 $Y=112830 $D=8
M1113 4805 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=399575 $Y=160970 $D=8
M1114 4806 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=399575 $Y=164845 $D=8
M1115 VDD 4630 4632 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=179690 $D=8
M1116 VDD 5306 5307 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=180970 $D=8
M1117 VDD 5314 5315 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=215690 $D=8
M1118 VDD 5370 5371 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=216970 $D=8
M1119 VDD 5378 5379 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=251690 $D=8
M1120 VDD 5478 5479 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=252970 $D=8
M1121 4630 4632 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=179690 $D=8
M1122 5306 5307 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=180970 $D=8
M1123 5314 5315 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=215690 $D=8
M1124 5370 5371 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=216970 $D=8
M1125 5378 5379 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=251690 $D=8
M1126 5478 5479 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=252970 $D=8
M1127 VDD 4466 4468 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=179690 $D=8
M1128 VDD 5328 5329 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=180970 $D=8
M1129 VDD 5336 5337 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=215690 $D=8
M1130 VDD 5392 5393 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=216970 $D=8
M1131 VDD 5400 5401 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=251690 $D=8
M1132 VDD 5492 5493 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=252970 $D=8
M1133 4786 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=402665 $Y=160970 $D=8
M1134 4785 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=402665 $Y=164845 $D=8
M1135 5426 4670 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=402880 $Y=112830 $D=8
M1136 4466 4468 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=179690 $D=8
M1137 5328 5329 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=180970 $D=8
M1138 5336 5337 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=215690 $D=8
M1139 5392 5393 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=216970 $D=8
M1140 5400 5401 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=251690 $D=8
M1141 5492 5493 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=252970 $D=8
M1142 5425 4671 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=405410 $Y=112830 $D=8
M1143 VDD 4462 4464 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=179690 $D=8
M1144 VDD 5326 5327 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=180970 $D=8
M1145 VDD 5334 5335 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=215690 $D=8
M1146 VDD 5390 5391 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=216970 $D=8
M1147 VDD 5398 5399 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=251690 $D=8
M1148 VDD 5490 5491 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=252970 $D=8
M1149 4783 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=405765 $Y=160970 $D=8
M1150 4784 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=405765 $Y=164845 $D=8
M1151 4462 4464 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=179690 $D=8
M1152 5326 5327 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=180970 $D=8
M1153 5334 5335 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=215690 $D=8
M1154 5390 5391 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=216970 $D=8
M1155 5398 5399 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=251690 $D=8
M1156 5490 5491 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=252970 $D=8
M1157 VDD 4458 4460 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=179690 $D=8
M1158 VDD 5324 5325 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=180970 $D=8
M1159 VDD 5332 5333 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=215690 $D=8
M1160 VDD 5388 5389 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=216970 $D=8
M1161 VDD 5396 5397 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=251690 $D=8
M1162 VDD 5488 5489 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=252970 $D=8
M1163 4782 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=408860 $Y=160970 $D=8
M1164 4781 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=408860 $Y=164845 $D=8
M1165 5424 4672 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=409075 $Y=112830 $D=8
M1166 4458 4460 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=179690 $D=8
M1167 5324 5325 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=180970 $D=8
M1168 5332 5333 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=215690 $D=8
M1169 5388 5389 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=216970 $D=8
M1170 5396 5397 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=251690 $D=8
M1171 5488 5489 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=252970 $D=8
M1172 VDD 4454 4456 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=179690 $D=8
M1173 VDD 5322 5323 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=180970 $D=8
M1174 VDD 5330 5331 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=215690 $D=8
M1175 VDD 5386 5387 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=216970 $D=8
M1176 VDD 5394 5395 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=251690 $D=8
M1177 VDD 5486 5487 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=252970 $D=8
M1178 5423 4673 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=411605 $Y=112830 $D=8
M1179 4779 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=411960 $Y=160970 $D=8
M1180 4780 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=411960 $Y=164845 $D=8
M1181 4454 4456 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=179690 $D=8
M1182 5322 5323 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=180970 $D=8
M1183 5330 5331 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=215690 $D=8
M1184 5386 5387 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=216970 $D=8
M1185 5394 5395 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=251690 $D=8
M1186 5486 5487 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=252970 $D=8
M1187 VDD VSS VDD VDD pfet_05v0 L=2.365e-06 W=8.19e-05 AD=0 AS=6.1309e-11 PD=0 PS=0.000217698 NRD=0 NRS=11.8457 m=1 nf=36 $X=304360 $Y=171065 $D=8
M1188 614 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=6.35965e-12 PD=7.86e-06 PS=1.737e-05 NRD=0.152493 NRS=0.546921 m=1 nf=2 $X=418655 $Y=160970 $D=8
M1189 615 936 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=6.35965e-12 PD=7.86e-06 PS=1.737e-05 NRD=0.152493 NRS=0.546921 m=1 nf=2 $X=418655 $Y=164845 $D=8
M1190 606 614 VDD VDD pfet_05v0 L=6e-07 W=7.02e-06 AD=1.8252e-12 AS=3.0888e-12 PD=8.06e-06 PS=1.58e-05 NRD=0.148148 NRS=0.250712 m=1 nf=2 $X=418770 $Y=97440 $D=8
M1191 607 606 VDD VDD pfet_05v0 L=6e-07 W=2.128e-05 AD=5.5328e-12 AS=9.3632e-12 PD=2.232e-05 PS=4.432e-05 NRD=0.0488722 NRS=0.0827068 m=1 nf=2 $X=418790 $Y=67070 $D=8
M1192 613 VDD VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=2.33887e-12 PD=4.29e-06 PS=9.09e-06 NRD=0.444444 NRS=1.06061 m=1 nf=2 $X=418870 $Y=112830 $D=8
X1198 614 614 613 VDD pfet_05v0_I04 $T=419815 124190 0 180 $X=418175 $Y=116760
X1199 615 615 613 VDD pfet_05v0_I04 $T=419815 151940 0 180 $X=418175 $Y=144510
X1200 615 614 936 VDD pfet_05v0_I04 $T=419825 159875 0 180 $X=418185 $Y=152445
X1201 614 614 VDD VSS nfet_05v0_I04 $T=419815 133465 0 180 $X=418535 $Y=126035
X1202 615 615 VDD VSS nfet_05v0_I04 $T=419815 143485 0 180 $X=418535 $Y=136055
X1208 VDD 618 616 pmos_1p2$$46273580 $T=242390 65835 1 0 $X=240960 $Y=64015
X1209 VSS 617 787 VSS nmos_1p2$$46563372 $T=233925 66830 0 0 $X=232780 $Y=66145
X1210 618 VSS 616 VSS nmos_1p2$$46563372 $T=243510 68190 1 0 $X=242365 $Y=66555
X1211 619 618 617 VSS nmos_1p2$$46563372 $T=246080 68190 1 0 $X=244935 $Y=66555
X1213 937 VSS Q[0] D[0] 4218 1 VDD 938 939 WEN[0] 4699 4700 4701 4702 4703 4704 4705 4706 4707 4708
+ 4709 4710 4711 4712 4818 927 4664 4663 4662 4661 4660 4659 4658 4657 4665 4862 4863 4864 4865 4866
+ 4867 4868
+ saout_m2 $T=9775 25090 0 0 $X=8430 $Y=7315
X1214 912 VSS Q[2] D[2] 4219 1 VDD 940 941 WEN[2] 4713 4714 4715 4716 4717 4718 4719 4720 4721 4722
+ 4723 4724 4725 4726 4819 927 4664 4663 4662 4661 4660 4659 4658 4657 4665 4869 4870 4871 4872 4873
+ 4874 4875
+ saout_m2 $T=63775 25090 0 0 $X=62430 $Y=7315
X1215 942 VSS Q[4] D[4] 4220 1 VDD 943 944 WEN[4] 4727 4728 4729 4730 4731 4732 4733 4734 4735 4736
+ 4737 4738 4739 4740 4820 927 4666 4667 4668 4669 4670 4671 4672 4673 4665 4876 4877 4878 4879 4880
+ 4881 4882
+ saout_m2 $T=307655 25090 0 0 $X=306310 $Y=7315
X1216 945 VSS Q[6] D[6] 4221 1 VDD 946 947 WEN[6] 4741 4742 4743 4744 4745 4746 4747 4748 4749 4750
+ 4751 4752 4753 4754 4821 927 4666 4667 4668 4669 4670 4671 4672 4673 4665 4883 4884 4885 4886 4887
+ 4888 4889
+ saout_m2 $T=361655 25090 0 0 $X=360310 $Y=7315
X1217 VSS VSS 4261 4262 4263 4264 4265 4266 4267 4268 ICV_4 $T=27210 176130 1 180 $X=23870 $Y=175790
X1218 VSS VSS 4269 4270 4271 4272 4273 4274 4275 4276 ICV_4 $T=33210 176130 1 180 $X=29870 $Y=175790
X1219 VSS VSS 4277 4278 4279 4280 4281 4282 4283 4284 ICV_4 $T=81210 176130 1 180 $X=77870 $Y=175790
X1220 VSS VSS 4285 4286 4287 4288 4289 4290 4291 4292 ICV_4 $T=87210 176130 1 180 $X=83870 $Y=175790
X1221 VSS VSS 4293 4294 4295 4296 4297 4298 4299 4300 ICV_4 $T=325090 176130 1 180 $X=321750 $Y=175790
X1222 VSS VSS 4301 4302 4303 4304 4305 4306 4307 4308 ICV_4 $T=331090 176130 1 180 $X=327750 $Y=175790
X1223 VSS VSS 4309 4310 4311 4312 4313 4314 4315 4316 ICV_4 $T=379090 176130 1 180 $X=375750 $Y=175790
X1224 VSS VSS 4317 4318 4319 4320 4321 4322 4323 4324 ICV_4 $T=385090 176130 1 180 $X=381750 $Y=175790
X1225 VSS VSS 4325 4326 4327 4328 4329 4330 4331 4332 4333 4334 4335 4336 4337 4338 4339 4340 ICV_5 $T=27210 257130 0 180 $X=23870 $Y=252290
X1226 VSS VSS 4341 4342 4343 4344 4345 4346 4347 4348 4349 4350 4351 4352 4353 4354 4355 4356 ICV_5 $T=54210 176130 1 180 $X=50870 $Y=175790
X1227 VSS VSS 4357 4358 4359 4360 4361 4362 4363 4364 4365 4366 4367 4368 4369 4370 4371 4372 ICV_5 $T=54210 257130 0 180 $X=50870 $Y=252290
X1228 VSS VSS 4373 4374 4375 4376 4377 4378 4379 4380 4381 4382 4383 4384 4385 4386 4387 4388 ICV_5 $T=108210 176130 1 180 $X=104870 $Y=175790
X1229 VSS 861 4389 4390 4391 4392 4393 4394 4395 4396 4397 4398 4399 4400 4401 4402 4403 4404 ICV_5 $T=313090 257130 0 180 $X=309750 $Y=252290
X1230 VSS 861 4405 4406 4407 4408 4409 4410 4411 4412 4413 4414 4415 4416 4417 4418 4419 4420 ICV_5 $T=325090 257130 0 180 $X=321750 $Y=252290
X1231 VSS VSS 4421 4422 4423 4424 4425 4426 4427 4428 4429 4430 4431 4432 4433 4434 4435 4436 ICV_5 $T=352090 176130 1 180 $X=348750 $Y=175790
X1232 VSS 861 4437 4438 4439 4440 4441 4442 4443 4444 4445 4446 4447 4448 4449 4450 4451 4452 ICV_5 $T=352090 257130 0 180 $X=348750 $Y=252290
X1233 VSS VSS 4453 4454 4455 4456 4457 4458 4459 4460 4461 4462 4463 4464 4465 4466 4467 4468 ICV_5 $T=406090 176130 1 180 $X=402750 $Y=175790
X1237 VSS VSS 4469 4470 4471 4472 4473 4474 4475 4476 4477 4478 4479 4480 4481 4482 4483 4484 ICV_7 $T=12210 176130 1 180 $X=8870 $Y=175790
X1238 VSS VSS 4485 4486 4487 4488 4489 4490 4491 4492 4493 4494 4495 4496 4497 4498 4499 4500 ICV_7 $T=12210 257130 0 180 $X=8870 $Y=252290
X1239 VSS VSS 4501 4502 4503 4504 4505 4506 4507 4508 4509 4510 4511 4512 4513 4514 4515 4516 ICV_7 $T=39210 176130 1 180 $X=35870 $Y=175790
X1240 VSS VSS 4517 4518 4519 4520 4521 4522 4523 4524 4525 4526 4527 4528 4529 4530 4531 4532 ICV_7 $T=39210 257130 0 180 $X=35870 $Y=252290
X1241 VSS VSS 4533 4534 4535 4536 4537 4538 4539 4540 4541 4542 4543 4544 4545 4546 4547 4548 ICV_7 $T=66210 176130 1 180 $X=62870 $Y=175790
X1242 VSS VSS 4549 4550 4551 4552 4553 4554 4555 4556 4557 4558 4559 4560 4561 4562 4563 4564 ICV_7 $T=93210 176130 1 180 $X=89870 $Y=175790
X1243 VSS VSS 4565 4566 4567 4568 4569 4570 4571 4572 4573 4574 4575 4576 4577 4578 4579 4580 ICV_7 $T=310090 176130 1 180 $X=306750 $Y=175790
X1244 VSS VSS 4581 4582 4583 4584 4585 4586 4587 4588 4589 4590 4591 4592 4593 4594 4595 4596 ICV_7 $T=337090 176130 1 180 $X=333750 $Y=175790
X1245 VSS 861 4597 4598 4599 4600 4601 4602 4603 4604 4605 4606 4607 4608 4609 4610 4611 4612 ICV_7 $T=337090 257130 0 180 $X=333750 $Y=252290
X1246 VSS VSS 4613 4614 4615 4616 4617 4618 4619 4620 4621 4622 4623 4624 4625 4626 4627 4628 ICV_7 $T=364090 176130 1 180 $X=360750 $Y=175790
X1247 VSS VSS 4629 4630 4631 4632 4633 4634 4635 4636 4637 4638 4639 4640 4641 4642 4643 4644 ICV_7 $T=391090 176130 1 180 $X=387750 $Y=175790
X1281 VDD VSS 4222 4223 4224 4225 4226 4227 4228 4229 4699 4700 4701 4702 4703 4704 4705 4706 4707 4708
+ 4709 4710 4711 4712 939 938 4787 4788 4789 4790 4791 4792 951 950 4755 4756 4757 4758 4759 4760
+ 4761 4762 4890 4891 4892 4893 4894 4895 4896 4897 4898 4899 4900 4901 4902 4903 4904 4905 4906 4907
+ 4908 4909 4910 4911 4912 4913 4914 4915 4916 4917 4918 4919 4920 4921 4922 4923 4924 4925 4926 4927
+ 4928 4929 4930 4931 4932 4933 4934 4935 4936 4937 4938 4939 4940 4941 4942 4943 4944 4945 4946 4947
+ 4948 4949 4950 4951 4952 4953
+ ICV_18 $T=12210 180630 0 0 $X=11870 $Y=180290
X1282 VDD VSS 4230 4231 4232 4233 4234 4235 4236 4237 4699 4700 4701 4702 4703 4704 4705 4706 4707 4708
+ 4709 4710 4711 4712 939 938 4787 4788 4789 4790 4791 4792 951 950 4755 4756 4757 4758 4759 4760
+ 4761 4762 4954 4955 4956 4957 4958 4959 4960 4961 4962 4963 4964 4965 4966 4967 4968 4969 4970 4971
+ 4972 4973 4974 4975 4976 4977 4978 4979 4980 4981 4982 4983 4984 4985 4986 4987 4988 4989 4990 4991
+ 4992 4993 4994 4995 4996 4997 4998 4999 5000 5001 5002 5003 5004 5005 5006 5007 5008 5009 5010 5011
+ 5012 5013 5014 5015 5016 5017
+ ICV_18 $T=12210 216630 0 0 $X=11870 $Y=216290
X1283 VDD VSS 4222 4223 4224 4225 4226 4227 4228 4229 4713 4714 4715 4716 4717 4718 4719 4720 4721 4722
+ 4723 4724 4725 4726 941 940 4793 4794 4795 4796 4797 4798 954 953 4763 4764 4765 4766 4767 4768
+ 4769 4770 5018 5019 5020 5021 5022 5023 5024 5025 5026 5027 5028 5029 5030 5031 5032 5033 5034 5035
+ 5036 5037 5038 5039 5040 5041 5042 5043 5044 5045 5046 5047 5048 5049 5050 5051 5052 5053 5054 5055
+ 5056 5057 5058 5059 5060 5061 5062 5063 5064 5065 5066 5067 5068 5069 5070 5071 5072 5073 5074 5075
+ 5076 5077 5078 5079 5080 5081
+ ICV_18 $T=66210 180630 0 0 $X=65870 $Y=180290
X1284 VDD VSS 4230 4231 4232 4233 4234 4235 4236 4237 4713 4714 4715 4716 4717 4718 4719 4720 4721 4722
+ 4723 4724 4725 4726 941 940 4793 4794 4795 4796 4797 4798 954 953 4763 4764 4765 4766 4767 4768
+ 4769 4770 5082 5083 5084 5085 5086 5087 5088 5089 5090 5091 5092 5093 5094 5095 5096 5097 5098 5099
+ 5100 5101 5102 5103 5104 5105 5106 5107 5108 5109 5110 5111 5112 5113 5114 5115 5116 5117 5118 5119
+ 5120 5121 5122 5123 5124 5125 5126 5127 5128 5129 5130 5131 5132 5133 5134 5135 5136 5137 5138 5139
+ 5140 5141 5142 5143 5144 5145
+ ICV_18 $T=66210 216630 0 0 $X=65870 $Y=216290
X1285 VDD VSS 4238 4239 4240 4241 4242 4243 4244 4245 4727 4728 4729 4730 4731 4732 4733 4734 4735 4736
+ 4737 4738 4739 4740 944 943 4799 4800 4801 4802 4803 4804 958 957 4771 4772 4773 4774 4775 4776
+ 4777 4778 5146 5147 5148 5149 5150 5151 5152 5153 5154 5155 5156 5157 5158 5159 5160 5161 5162 5163
+ 5164 5165 5166 5167 5168 5169 5170 5171 5172 5173 5174 5175 5176 5177 5178 5179 5180 5181 5182 5183
+ 5184 5185 5186 5187 5188 5189 5190 5191 5192 5193 5194 5195 5196 5197 5198 5199 5200 5201 5202 5203
+ 5204 5205 5206 5207 5208 5209
+ ICV_18 $T=310090 180630 0 0 $X=309750 $Y=180290
X1286 VDD VSS 4246 4247 4248 4249 4250 4251 4252 4253 4727 4728 4729 4730 4731 4732 4733 4734 4735 4736
+ 4737 4738 4739 4740 944 943 4799 4800 4801 4802 4803 4804 958 957 4771 4772 4773 4774 4775 4776
+ 4777 4778 5210 5211 5212 5213 5214 5215 5216 5217 5218 5219 5220 5221 5222 5223 5224 5225 5226 5227
+ 5228 5229 5230 5231 5232 5233 5234 5235 5236 5237 5238 5239 5240 5241 5242 5243 5244 5245 5246 5247
+ 5248 5249 5250 5251 5252 5253 5254 5255 5256 5257 5258 5259 5260 5261 5262 5263 5264 5265 5266 5267
+ 5268 5269 5270 5271 5272 5273
+ ICV_18 $T=310090 216630 0 0 $X=309750 $Y=216290
X1287 VDD VSS 4238 4239 4240 4241 4242 4243 4244 4245 4741 4742 4743 4744 4745 4746 4747 4748 4749 4750
+ 4751 4752 4753 4754 947 946 4805 4806 4807 4808 4809 4810 961 960 4779 4780 4781 4782 4783 4784
+ 4785 4786 5274 5275 5276 5277 5278 5279 5280 5281 5282 5283 5284 5285 5286 5287 5288 5289 5290 5291
+ 5292 5293 5294 5295 5296 5297 5298 5299 5300 5301 5302 5303 5304 5305 5306 5307 5308 5309 5310 5311
+ 5312 5313 5314 5315 5316 5317 5318 5319 5320 5321 5322 5323 5324 5325 5326 5327 5328 5329 5330 5331
+ 5332 5333 5334 5335 5336 5337
+ ICV_18 $T=364090 180630 0 0 $X=363750 $Y=180290
X1288 VDD VSS 4246 4247 4248 4249 4250 4251 4252 4253 4741 4742 4743 4744 4745 4746 4747 4748 4749 4750
+ 4751 4752 4753 4754 947 946 4805 4806 4807 4808 4809 4810 961 960 4779 4780 4781 4782 4783 4784
+ 4785 4786 5338 5339 5340 5341 5342 5343 5344 5345 5346 5347 5348 5349 5350 5351 5352 5353 5354 5355
+ 5356 5357 5358 5359 5360 5361 5362 5363 5364 5365 5366 5367 5368 5369 5370 5371 5372 5373 5374 5375
+ 5376 5377 5378 5379 5380 5381 5382 5383 5384 5385 5386 5387 5388 5389 5390 5391 5392 5393 5394 5395
+ 5396 5397 5398 5399 5400 5401
+ ICV_18 $T=364090 216630 0 0 $X=363750 $Y=216290
X1289 949 VSS Q[1] 948 D[1] 1 VDD 950 951 WEN[1] 4755 4756 4757 4758 4759 4760 4761 4762 4787 4788
+ 4789 4790 4791 4792 4822 4657 4658 4659 927 4660 4661 4662 4663 4664 4665 5402 5403 5404 5405 5406
+ 5407 5408
+ saout_R_m2 $T=65645 25125 1 180 $X=27480 $Y=6815
X1290 913 VSS Q[3] 952 D[3] 1 VDD 953 954 WEN[3] 4763 4764 4765 4766 4767 4768 4769 4770 4793 4794
+ 4795 4796 4797 4798 4823 4657 4658 4659 927 4660 4661 4662 4663 4664 4665 5409 5410 5411 5412 5413
+ 5414 5415
+ saout_R_m2 $T=119645 25125 1 180 $X=81480 $Y=6815
X1291 956 VSS Q[5] 955 D[5] 1 VDD 957 958 WEN[5] 4771 4772 4773 4774 4775 4776 4777 4778 4799 4800
+ 4801 4802 4803 4804 4824 4673 4672 4671 927 4670 4669 4668 4667 4666 4665 5416 5417 5418 5419 5420
+ 5421 5422
+ saout_R_m2 $T=363525 25125 1 180 $X=325360 $Y=6815
X1292 959 VSS Q[7] 936 D[7] 1 VDD 960 961 WEN[7] 4779 4780 4781 4782 4783 4784 4785 4786 4805 4806
+ 4807 4808 4809 4810 4825 4673 4672 4671 927 4670 4669 4668 4667 4666 4665 5423 5424 5425 5426 5427
+ 5428 5429
+ saout_R_m2 $T=417525 25125 1 180 $X=379360 $Y=6815
X1293 VSS VSS 5430 5431 5432 5433 5434 5435 5436 5437 5438 5439 5440 5441 5442 5443 5444 5445 5446 5447
+ 5448 5449 5450 5451 5452 5453 5454 5455 5456 5457 5458 5459 5460 5461
+ new_dummyrow_unit $T=65900 258015 1 0 $X=65870 $Y=252290
X1294 VSS 861 5462 5463 5464 5465 5466 5467 5468 5469 5470 5471 5472 5473 5474 5475 5476 5477 5478 5479
+ 5480 5481 5482 5483 5484 5485 5486 5487 5488 5489 5490 5491 5492 5493
+ new_dummyrow_unit $T=363780 258015 1 0 $X=363750 $Y=252290
X1297 732 733 VSS 5494 5495 5496 5497 ICV_24 $T=117210 185130 0 0 $X=116870 $Y=180290
X1298 732 733 VSS 5498 5499 5500 5501 ICV_24 $T=117210 194130 0 0 $X=116870 $Y=189290
X1299 732 733 VSS 5502 5503 5504 5505 ICV_24 $T=117210 203130 0 0 $X=116870 $Y=198290
X1300 732 733 VSS 5506 5507 5508 5509 ICV_24 $T=117210 212130 0 0 $X=116870 $Y=207290
X1301 732 733 VSS 5510 5511 5512 5513 ICV_24 $T=117210 221130 0 0 $X=116870 $Y=216290
X1302 732 733 VSS 5514 5515 5516 5517 ICV_24 $T=117210 230130 0 0 $X=116870 $Y=225290
X1303 732 733 VSS 5518 5519 5520 5521 ICV_24 $T=117210 239130 0 0 $X=116870 $Y=234290
X1304 732 733 VSS 5522 5523 5524 5525 ICV_24 $T=117210 248130 0 0 $X=116870 $Y=243290
X1322 VSS VDD 1 CLK VSS VSS 4682 4683 4687 4688 xpredec0 $T=146075 111460 0 0 $X=144630 $Y=111455
X1323 VSS VDD 1 CLK VSS A[6] 4689 4690 917 918 xpredec0 $T=182970 111460 0 0 $X=181525 $Y=111455
X1328 VSS VDD 1 CLK 4663 4664 4657 4658 4659 4660 4661 4662 4673 4672 4671 4670 4669 4668 4667 4666
+ A[2] A[1] A[0]
+ ypredec1 $T=145470 26355 0 0 $X=146365 $Y=26735
X1329 VSS VDD 918 925 924 923 922 921 920 VDD 4826 1 4827 4223 4239 4224 4240 4225 4241 4226
+ 4242 4227 4243 4228 4244 4828 4829 4854 4855 4856 4857
+ xdec8 $T=152015 180635 0 0 $X=152015 $Y=179495
X1330 VSS VDD 917 925 924 923 922 921 920 VDD 4830 1 4831 4231 4247 4232 4248 4233 4249 4234
+ 4250 4235 4251 4236 4252 4832 4833 4858 4859 4860 4861
+ xdec8 $T=152015 216635 0 0 $X=152015 $Y=215495
X1333 860 VSS 862 nfet_05v0_I19 $T=175115 254995 0 90 $X=164385 $Y=254315
X1334 861 VSS 863 nfet_05v0_I19 $T=260115 254995 0 90 $X=249385 $Y=254315
X1338 VDD 860 862 pmos_1p2$$204216364 $T=189610 255150 0 90 $X=176320 $Y=253670
X1339 VDD 861 863 pmos_1p2$$204216364 $T=248135 255150 0 90 $X=234845 $Y=253670
X1340 862 VDD 2 VDD pfet_05v0_I17 $T=198405 254995 0 90 $X=191195 $Y=253955
X1341 1 2 VSS VDD pfet_05v0_I17 $T=219905 254995 0 90 $X=212695 $Y=253955
X1342 863 VDD 2 VDD pfet_05v0_I17 $T=233255 254995 0 90 $X=226045 $Y=253955
X1343 862 VSS 2 nfet_05v0_I09 $T=202950 254995 0 90 $X=199690 $Y=254315
X1344 863 VSS 2 nfet_05v0_I09 $T=224800 254995 0 90 $X=221540 $Y=254315
X1345 VSS VDD GWEN CLK 4665 927 wen_v2 $T=208415 16605 0 0 $X=208280 $Y=15275
X1346 VSS 1 VDD CLK A[5] A[4] A[3] 919 920 921 922 923 924 925 926 xpredec1 $T=219860 111460 0 0 $X=219855 $Y=111455
X1347 VDD 864 CLK pfet_05v0_I06 $T=234280 43425 1 0 $X=233240 $Y=41905
X1348 VDD 865 864 pfet_05v0_I06 $T=239670 43425 1 0 $X=238630 $Y=41905
X1349 VSS 864 CLK nfet_05v0_I10 $T=234280 46585 1 0 $X=233600 $Y=45365
X1350 VSS 865 864 nfet_05v0_I10 $T=239670 46585 1 0 $X=238990 $Y=45365
X1370 VSS 734 735 5534 5535 5536 5537 ICV_19 $T=307090 180630 1 180 $X=303750 $Y=180290
X1371 VSS 734 735 5538 5539 5540 5541 ICV_19 $T=307090 189630 1 180 $X=303750 $Y=189290
X1372 VSS 734 735 5542 5543 5544 5545 ICV_19 $T=307090 198630 1 180 $X=303750 $Y=198290
X1373 VSS 734 735 5546 5547 5548 5549 ICV_19 $T=307090 207630 1 180 $X=303750 $Y=207290
X1374 VSS 734 735 5550 5551 5552 5553 ICV_19 $T=307090 216630 1 180 $X=303750 $Y=216290
X1375 VSS 734 735 5554 5555 5556 5557 ICV_19 $T=307090 225630 1 180 $X=303750 $Y=225290
X1376 VSS 734 735 5558 5559 5560 5561 ICV_19 $T=307090 234630 1 180 $X=303750 $Y=234290
X1377 VSS 734 735 5562 5563 5564 5565 ICV_19 $T=307090 243630 1 180 $X=303750 $Y=243290
X1379 VSS VDD 4834 4835 4836 4837 ICV_1 $T=418090 248130 0 0 $X=417750 $Y=247790
X1380 614 615 VSS VDD 4838 4839 4840 4841 ICV_2 $T=418090 176130 0 0 $X=417750 $Y=175790
X1381 614 615 VSS VDD 4842 4843 4844 4845 ICV_2 $T=418090 194130 0 0 $X=417750 $Y=193790
X1382 614 615 VSS VDD 4846 4847 4848 4849 ICV_2 $T=418090 212130 0 0 $X=417750 $Y=211790
X1383 614 615 VSS VDD 4850 4851 4852 4853 ICV_2 $T=418090 230130 0 0 $X=417750 $Y=229790
.ENDS
