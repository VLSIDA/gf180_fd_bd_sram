* Subcircuit definition of cell ICV_15
.SUBCKT ICV_15 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36 37
** N=53 EP=33 IP=55 FDC=32
*.SEEDPROM
X0 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 ICV_13 $T=-15000 0 0 0 $X=-24340 $Y=-340
X1 4 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 ICV_14 $T=0 0 0 0 $X=-12340 $Y=-340
.ENDS
