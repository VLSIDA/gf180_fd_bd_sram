* Subcircuit definition of cell 018SRAM_strap1_2x
.SUBCKT 018SRAM_strap1_2x
** N=10 EP=0 IP=12 FDC=0
.ENDS
