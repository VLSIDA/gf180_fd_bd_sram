* Subcircuit definition of cell ICV_28
.SUBCKT ICV_28 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=26 EP=18 IP=32 FDC=40
*.SEEDPROM
M0 1 20 19 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=8060 $D=8
M1 1 24 23 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=9340 $D=8
M2 20 19 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=8060 $D=8
M3 24 23 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=9340 $D=8
M4 1 22 21 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=8060 $D=8
M5 1 26 25 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=9340 $D=8
M6 22 21 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=8060 $D=8
M7 26 25 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=9340 $D=8
X8 2 3 4 7 8 9 10 11 19 12 20 13 21 14 22 ICV_27 $T=0 0 0 0 $X=-340 $Y=-340
X9 2 5 6 7 8 9 10 23 15 24 16 25 17 26 18 ICV_27 $T=0 9000 0 0 $X=-340 $Y=8660
.ENDS
