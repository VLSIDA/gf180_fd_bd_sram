* Subcircuit definition of cell ICV_22
.SUBCKT ICV_22 1 2 5 8 9 10 11 12
** N=22 EP=8 IP=36 FDC=16
M0 20 10 13 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=1.73655e-12 AS=4.05195e-12 PD=7.32e-06 PS=1.481e-05 NRD=0.0374449 NRS=0.0873715 m=1 nf=1 $X=-2370 $Y=-33035 $D=2
M1 19 9 20 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=3.405e-14 AS=-3.405e-14 PD=1e-08 PS=-1e-08 NRD=0.000734214 NRS=-0.000734214 m=1 nf=1 $X=-1260 $Y=-33035 $D=2
M2 1 2 19 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=3.405e-14 AS=-3.405e-14 PD=1e-08 PS=-1e-08 NRD=0.000734214 NRS=-0.000734214 m=1 nf=1 $X=-140 $Y=-33035 $D=2
M3 1 13 11 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=1.7706e-12 AS=2.1792e-12 PD=8.37e-06 PS=1.1e-05 NRD=0.343612 NRS=0.422907 m=1 nf=3 $X=-2375 $Y=-2950 $D=2
M4 21 5 1 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=-3.405e-14 AS=3.405e-14 PD=-1e-08 PS=1e-08 NRD=-0.000734214 NRS=0.000734214 m=1 nf=1 $X=990 $Y=-33035 $D=2
M5 22 9 21 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=-3.405e-14 AS=3.405e-14 PD=-1e-08 PS=1e-08 NRD=-0.000734214 NRS=0.000734214 m=1 nf=1 $X=2110 $Y=-33035 $D=2
M6 16 10 22 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=4.05195e-12 AS=1.73655e-12 PD=1.481e-05 PS=7.32e-06 NRD=0.0873715 NRS=0.0374449 m=1 nf=1 $X=3220 $Y=-33035 $D=2
M7 12 16 1 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=2.1792e-12 AS=1.7706e-12 PD=1.1e-05 PS=8.37e-06 NRD=0.422907 NRS=0.343612 m=1 nf=3 $X=985 $Y=-2950 $D=2
M8 8 10 13 8 pfet_05v0 L=6e-07 W=5.67e-06 AD=1.4742e-12 AS=2.4948e-12 PD=6.19e-06 PS=1.222e-05 NRD=0.0458554 NRS=0.0776014 m=1 nf=1 $X=-2375 $Y=-19360 $D=8
M9 13 9 8 8 pfet_05v0 L=6e-07 W=5.67e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=-1255 $Y=-19360 $D=8
M10 8 2 13 8 pfet_05v0 L=6e-07 W=5.67e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=-135 $Y=-19360 $D=8
M11 8 13 11 8 pfet_05v0 L=6e-07 W=1.731e-05 AD=4.5006e-12 AS=5.5392e-12 PD=1.887e-05 PS=2.5e-05 NRD=0.135182 NRS=0.166378 m=1 nf=3 $X=-2375 $Y=-10125 $D=8
M12 16 5 8 8 pfet_05v0 L=6e-07 W=5.67e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=985 $Y=-19360 $D=8
M13 8 9 16 8 pfet_05v0 L=6e-07 W=5.67e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=2105 $Y=-19360 $D=8
M14 16 10 8 8 pfet_05v0 L=6e-07 W=5.67e-06 AD=2.4948e-12 AS=1.4742e-12 PD=1.222e-05 PS=6.19e-06 NRD=0.0776014 NRS=0.0458554 m=1 nf=1 $X=3225 $Y=-19360 $D=8
M15 12 16 8 8 pfet_05v0 L=6e-07 W=1.731e-05 AD=5.5392e-12 AS=4.5006e-12 PD=2.5e-05 PS=1.887e-05 NRD=0.166378 NRS=0.135182 m=1 nf=3 $X=985 $Y=-10125 $D=8
.ENDS
