* Subcircuit definition of cell xdec
.SUBCKT xdec 1 2 men 6 vss 8 28 vdd
** N=98 EP=8 IP=41 FDC=6
*.SEEDPROM
M0 2 6 men vss nfet_05v0 L=6e-07 W=6.6e-06 AD=2.904e-12 AS=1.716e-12 PD=1.496e-05 PS=7.64e-06 NRD=0.266667 NRS=0.157576 m=1 nf=2 $X=37460 $Y=965 $D=2
M1 vss 8 6 vss nfet_05v0 L=6e-07 W=6.6e-07 AD=2.904e-13 AS=2.904e-13 PD=2.2e-06 PS=2.2e-06 NRD=0.666667 NRS=0.666667 m=1 nf=1 $X=45970 $Y=965 $D=2
M2 2 8 men vdd pfet_05v0 L=6e-07 W=6.6e-06 AD=2.904e-12 AS=1.716e-12 PD=1.496e-05 PS=7.64e-06 NRD=0.266667 NRS=0.157576 m=1 nf=2 $X=32185 $Y=965 $D=8
M3 vdd 8 6 vdd pfet_05v0 L=6e-07 W=1.59e-06 AD=6.996e-13 AS=6.996e-13 PD=4.06e-06 PS=4.06e-06 NRD=0.27673 NRS=0.27673 m=1 nf=1 $X=43020 $Y=965 $D=8
X12 vdd 1 2 pmos_1p2$$49272876_R270 $T=29780 1120 0 90 $X=23605 $Y=-360
X13 vdd 28 2 pmos_1p2$$49272876_R270 $T=91805 1120 1 90 $X=91120 $Y=-360
.ENDS
************* SUBCKT CALLS DEFINITION ***************
.SUBCKT pmos_1p2$$49272876_R270 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=1.1e-05 AD=2.86e-12 AS=4.84e-12 PD=1.204e-05 PS=2.376e-05 NRD=0.0945455 NRS=0.16 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
