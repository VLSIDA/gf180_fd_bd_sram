* Subcircuit definition of cell outbuf_oe
.SUBCKT outbuf_oe q vss 3 4 5 15 16 17 18 vdd GWE se qp qn 24
** N=66 EP=15 IP=48 FDC=18
M0 vss 5 q vss nfet_05v0 L=6e-07 W=1.272e-05 AD=3.3072e-12 AS=4.0704e-12 PD=1.584e-05 PS=2.08e-05 NRD=0.735849 NRS=0.90566 m=1 nf=6 $X=395 $Y=2665 $D=2
M1 3 GWE vss vss nfet_05v0 L=6e-07 W=1.6e-06 AD=7.04e-13 AS=7.04e-13 PD=4.08e-06 PS=4.08e-06 NRD=0.275 NRS=0.275 m=1 nf=1 $X=8145 $Y=2720 $D=2
M2 17 3 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=10105 $Y=2700 $D=2
M3 vss 16 4 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=13175 $Y=12845 $D=2
M4 5 15 4 vss nfet_05v0 L=6e-07 W=6.81e-06 AD=2.1792e-12 AS=2.1792e-12 PD=1.1e-05 PS=1.1e-05 NRD=0.422907 NRS=0.422907 m=1 nf=3 $X=12455 $Y=2720 $D=2
M5 vss se 15 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=17045 $Y=4035 $D=2
M6 5 qn 18 vss nfet_05v0 L=6e-07 W=5.68e-06 AD=1.4768e-12 AS=1.988e-12 PD=6.72e-06 PS=9.92e-06 NRD=0.183099 NRS=0.246479 m=1 nf=2 $X=19905 $Y=1945 $D=2
M7 vss 3 18 vss nfet_05v0 L=6e-07 W=5.68e-06 AD=1.4768e-12 AS=1.988e-12 PD=6.72e-06 PS=9.92e-06 NRD=0.183099 NRS=0.246479 m=1 nf=2 $X=22145 $Y=1945 $D=2
M8 vdd 5 q vdd pfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=7.2576e-12 PD=2.58e-05 PS=3.408e-05 NRD=0.412698 NRS=0.507937 m=1 nf=6 $X=395 $Y=6190 $D=8
M9 3 GWE vdd vdd pfet_05v0 L=6e-07 W=4e-06 AD=1.76e-12 AS=1.76e-12 PD=8.88e-06 PS=8.88e-06 NRD=0.11 NRS=0.11 m=1 nf=1 $X=8145 $Y=6395 $D=8
M10 17 3 vdd vdd pfet_05v0 L=6e-07 W=4.5e-06 AD=1.98e-12 AS=1.98e-12 PD=9.88e-06 PS=9.88e-06 NRD=0.0977778 NRS=0.0977778 m=1 nf=1 $X=10105 $Y=6175 $D=8
M11 4 16 vdd vdd pfet_05v0 L=6e-07 W=2.28e-06 AD=5.928e-13 AS=1.24202e-12 PD=3.32e-06 PS=5.60564e-06 NRD=0.45614 NRS=0.955691 m=1 nf=2 $X=12055 $Y=10310 $D=8
M12 5 se 4 vdd pfet_05v0 L=6e-07 W=6.81e-06 AD=2.1792e-12 AS=2.1792e-12 PD=1.1e-05 PS=1.1e-05 NRD=0.422907 NRS=0.422907 m=1 nf=3 $X=12455 $Y=6395 $D=8
M13 16 5 vdd vdd pfet_05v0 L=6e-07 W=1.2e-06 AD=5.28e-13 AS=7.79385e-13 PD=3.28e-06 PS=2.57436e-06 NRD=0.366667 NRS=0.541239 m=1 nf=1 $X=15085 $Y=10250 $D=8
M14 vdd se 15 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=17045 $Y=7030 $D=8
M15 5 qp 24 vdd pfet_05v0 L=6e-07 W=1.134e-05 AD=2.9484e-12 AS=3.969e-12 PD=1.238e-05 PS=1.841e-05 NRD=0.0917108 NRS=0.123457 m=1 nf=2 $X=19680 $Y=6685 $D=8
M16 vdd 17 24 vdd pfet_05v0 L=6e-07 W=1.134e-05 AD=2.9484e-12 AS=3.969e-12 PD=1.238e-05 PS=1.841e-05 NRD=0.0917108 NRS=0.123457 m=1 nf=2 $X=21920 $Y=6685 $D=8
X22 vss 16 5 vss nfet_05v0_I05 $T=15150 13365 1 0 $X=14470 $Y=12145
.ENDS
