* Subcircuit definition of cell ICV_37
.SUBCKT ICV_37 1 50 51 52 54 55 56 57 58 59 104 105 106 107 108 109 112 113 114 115
+ 116 117 119 126 127 128 129 130 131 132 133
** N=137 EP=31 IP=157 FDC=126
*.SEEDPROM
X0 1 51 52 59 58 57 56 55 54 50 126 119 127 104 112 105 113 106 114 107
+ 115 108 116 109 117 128 129 130 131 132 133
+ xdec8 $T=9750 2385 1 270 $X=-27390 $Y=-118710
.ENDS
