* Subcircuit definition of cell ICV_24
.SUBCKT ICV_24 1 50 94 95 96 100 101 114 117 118 121
** N=125 EP=11 IP=142 FDC=12
*.SEEDPROM
X0 114 94 95 115 1 96 117 50 xdec $T=0 0 1 0 $X=-5 $Y=-5640
X1 118 100 95 119 1 101 121 50 xdec $T=0 0 0 0 $X=-5 $Y=-1115
.ENDS
