* Subcircuit definition of cell 018SRAM_cell1
.SUBCKT 018SRAM_cell1
** N=8 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
