* Subcircuit definition of cell xpredec1_bot
.SUBCKT xpredec1_bot 1 2 3 10 11 12 13
** N=32 EP=7 IP=19 FDC=12
X0 1 32 11 10 13 12 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
X2 10 2 32 pmos_1p2$$47337516 $T=3910 18340 0 0 $X=2480 $Y=17635
X3 10 3 2 pmos_1p2$$47337516 $T=6480 18340 0 0 $X=5050 $Y=17635
X4 1 2 32 nmos_1p2$$47336492 $T=3910 36070 0 0 $X=2765 $Y=35385
X5 1 3 2 nmos_1p2$$47336492 $T=6480 36070 0 0 $X=5335 $Y=35385
.ENDS
************* SUBCKT CALLS DEFINITION ***************
.SUBCKT alatch vss ab a vdd enb en
** N=16 EP=6 IP=24 FDC=8
M0 ab 12 vss vss nfet_05v0 L=6e-07 W=3.64e-06 AD=9.464e-13 AS=1.6016e-12 PD=4.68e-06 PS=9.04e-06 NRD=0.285714 NRS=0.483516 m=1 nf=2 $X=2590 $Y=1475 $D=2
M1 vss ab 11 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=3710 $Y=12935 $D=2
M2 a en 12 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=6280 $Y=1020 $D=2
M3 11 enb 12 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=6280 $Y=12935 $D=2
M4 ab 12 vdd vdd pfet_05v0 L=6e-07 W=9.08e-06 AD=2.3608e-12 AS=3.9952e-12 PD=1.012e-05 PS=1.992e-05 NRD=0.114537 NRS=0.193833 m=1 nf=2 $X=2590 $Y=4695 $D=8
M5 a enb 12 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=6280 $Y=5895 $D=8
X10 11 vdd ab vdd pmos_1p2_161 $T=3865 11540 1 0 $X=2435 $Y=9910
X11 12 11 en vdd pmos_1p2_161 $T=6435 11540 1 0 $X=5005 $Y=9910
.ENDS
.SUBCKT pmos_1p2$$47337516 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=1.633e-05 AD=7.1852e-12 AS=7.1852e-12 PD=3.354e-05 PS=3.354e-05 NRD=0.0269443 NRS=0.0269443 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
.SUBCKT nmos_1p2$$47336492 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nfet_05v0 L=6e-07 W=6.58e-06 AD=2.8952e-12 AS=2.8952e-12 PD=1.404e-05 PS=1.404e-05 NRD=0.0668693 NRS=0.0668693 m=1 nf=1 $X=-155 $Y=0 $D=2
.ENDS
.SUBCKT pmos_1p2_161 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
M0 2 3 1 4 pfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
