* Subcircuit definition of cell sa
.SUBCKT sa 1 vss 3 4 qn qp 7 pcb vdd d db se
** N=105 EP=12 IP=47 FDC=27
M0 1 vss vss vss nfet_05v0 L=6e-07 W=3.41e-06 AD=8.866e-13 AS=1.5004e-12 PD=3.93e-06 PS=7.7e-06 NRD=0.0762463 NRS=0.129032 m=1 nf=1 $X=11660 $Y=16585 $D=2
M1 3 4 1 vss nfet_05v0 L=6e-07 W=3.41e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12780 $Y=16585 $D=2
M2 4 1 3 vss nfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=1.7732e-12 PD=7.86e-06 PS=7.86e-06 NRD=0.152493 NRS=0.152493 m=1 nf=2 $X=13900 $Y=16585 $D=2
M3 7 4 vss vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=15170 $Y=8510 $D=2
M4 1 4 3 vss nfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=1.7732e-12 PD=7.86e-06 PS=7.86e-06 NRD=0.152493 NRS=0.152493 m=1 nf=2 $X=16140 $Y=16585 $D=2
M5 4 1 3 vss nfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=1.7732e-12 PD=7.86e-06 PS=7.86e-06 NRD=0.152493 NRS=0.152493 m=1 nf=2 $X=18380 $Y=16585 $D=2
M6 vss 7 qp vss nfet_05v0 L=6e-07 W=6.81e-06 AD=1.7706e-12 AS=2.1792e-12 PD=8.37e-06 PS=1.1e-05 NRD=0.343612 NRS=0.422907 m=1 nf=3 $X=17410 $Y=8510 $D=2
M7 1 4 3 vss nfet_05v0 L=6e-07 W=3.41e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=20620 $Y=16585 $D=2
M8 qn 1 vss vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=20770 $Y=8510 $D=2
M9 3 se vss vss nfet_05v0 L=6e-07 W=2.272e-05 AD=5.9072e-12 AS=6.9296e-12 PD=2.688e-05 PS=3.328e-05 NRD=0.732394 NRS=0.859155 m=1 nf=8 $X=12945 $Y=12550 $D=2
M10 vss vss 1 vss nfet_05v0 L=6e-07 W=3.41e-06 AD=1.5004e-12 AS=8.866e-13 PD=7.7e-06 PS=3.93e-06 NRD=0.129032 NRS=0.0762463 m=1 nf=1 $X=21740 $Y=16585 $D=2
M11 4 vdd vdd vdd pfet_05v0 L=6e-07 W=9.1e-07 AD=2.366e-13 AS=4.004e-13 PD=1.43e-06 PS=2.7e-06 NRD=0.285714 NRS=0.483516 m=1 nf=1 $X=13985 $Y=24010 $D=8
M12 vdd 1 4 vdd pfet_05v0 L=6e-07 W=9.1e-07 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=15105 $Y=24010 $D=8
M13 d pcb vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=15755 $Y=30660 $D=8
M14 7 4 vdd vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.589e-12 PD=5.58e-06 PS=8.21e-06 NRD=0.229075 NRS=0.30837 m=1 nf=2 $X=15170 $Y=4385 $D=8
M15 4 pcb 1 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=16875 $Y=26330 $D=8
M16 db pcb d vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=16875 $Y=30660 $D=8
M17 1 4 vdd vdd pfet_05v0 L=6e-07 W=1.82e-06 AD=4.732e-13 AS=4.732e-13 PD=2.86e-06 PS=2.86e-06 NRD=0.571429 NRS=0.571429 m=1 nf=2 $X=16225 $Y=24010 $D=8
M18 vdd pcb db vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=17995 $Y=30660 $D=8
M19 4 1 vdd vdd pfet_05v0 L=6e-07 W=9.1e-07 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=18465 $Y=24010 $D=8
M20 qp 7 vdd vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.1804e-12 PD=5.58e-06 PS=5.58e-06 NRD=0.229075 NRS=0.229075 m=1 nf=2 $X=17410 $Y=4385 $D=8
M21 vdd vdd 4 vdd pfet_05v0 L=6e-07 W=9.1e-07 AD=4.004e-13 AS=2.366e-13 PD=2.7e-06 PS=1.43e-06 NRD=0.483516 NRS=0.285714 m=1 nf=1 $X=19585 $Y=24010 $D=8
M22 qn 1 vdd vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.589e-12 PD=5.58e-06 PS=8.21e-06 NRD=0.229075 NRS=0.30837 m=1 nf=2 $X=19650 $Y=4385 $D=8
X28 db 1 se vdd pmos_1p2$$46897196 $T=12475 26330 0 0 $X=11045 $Y=25620
X29 d 4 se vdd pmos_1p2$$46897196 $T=12475 30660 0 0 $X=11045 $Y=29950
X30 d 4 se vdd pmos_1p2$$46897196 $T=20400 26330 0 0 $X=18970 $Y=25620
X31 db 1 se vdd pmos_1p2$$46897196 $T=20400 30660 0 0 $X=18970 $Y=29950
.ENDS
************* SUBCKT CALLS DEFINITION ***************
.SUBCKT pmos_1p2$$46897196 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
M0 2 3 1 4 pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
