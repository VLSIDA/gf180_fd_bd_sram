* Subcircuit definition of cell ICV_41
.SUBCKT ICV_41 7 8 17 18 22 23 24 25
** N=29 EP=8 IP=48 FDC=44
*.SEEDPROM
M0 7 26 27 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=12560 $D=8
M1 7 28 29 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=13840 $D=8
M2 26 27 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=12560 $D=8
M3 28 29 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=13840 $D=8
X6 7 8 17 18 26 27 22 23 ICV_40 $T=6000 0 0 180 $X=2660 $Y=-4840
X7 7 8 17 18 24 25 28 29 ICV_40 $T=6000 18000 0 180 $X=2660 $Y=13160
.ENDS
