* Subcircuit definition of cell ICV_18
.SUBCKT ICV_18 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
** N=16 EP=15 IP=24 FDC=16
*.SEEDPROM
X0 5 6 2 3 4 9 11 10 12 018SRAM_cell1_2x $T=-3000 0 0 0 $X=-3340 $Y=-340
X1 7 8 2 3 4 13 15 14 16 018SRAM_cell1_2x $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
