* Subcircuit definition of cell nmos_1p2$$47514668
.SUBCKT nmos_1p2$$47514668
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
