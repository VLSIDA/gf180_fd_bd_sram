* Subcircuit definition of cell ypredec1
.SUBCKT ypredec1 1 2 men clk ly[6] ly[7] ly[0] ly[1] ly[2] ly[3] ly[4] ly[5] ry[0] ry[1] ry[2] ry[3] ry[4] ry[5] ry[6] ry[7]
+ A[2] A[1] A[0]
** N=374 EP=23 IP=151 FDC=172
M0 367 358 1 1 nfet_05v0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=3.9952e-12 PD=1.904e-05 PS=1.904e-05 NRD=0.0484581 NRS=0.0484581 m=1 nf=1 $X=2545 $Y=46970 $D=2
M1 1 371 ly[3] 1 nfet_05v0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=21585 $Y=46970 $D=2
M2 368 361 1 1 nfet_05v0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=24945 $Y=46970 $D=2
M3 188 189 1 1 nfet_05v0 L=6e-07 W=1.36e-06 AD=5.984e-13 AS=5.984e-13 PD=3.6e-06 PS=3.6e-06 NRD=0.323529 NRS=0.323529 m=1 nf=1 $X=31760 $Y=4985 $D=2
M4 189 clk 1 1 nfet_05v0 L=6e-07 W=1.91e-06 AD=4.966e-13 AS=8.404e-13 PD=2.43e-06 PS=4.7e-06 NRD=0.136126 NRS=0.230366 m=1 nf=1 $X=38610 $Y=5010 $D=2
M5 1 men 189 1 nfet_05v0 L=6e-07 W=1.91e-06 AD=8.404e-13 AS=4.966e-13 PD=4.7e-06 PS=2.43e-06 NRD=0.230366 NRS=0.136126 m=1 nf=1 $X=39730 $Y=5010 $D=2
M6 1 372 ly[7] 1 nfet_05v0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=43985 $Y=46970 $D=2
M7 369 358 1 1 nfet_05v0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=47345 $Y=46970 $D=2
M8 1 373 ry[3] 1 nfet_05v0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=66385 $Y=46970 $D=2
M9 370 361 1 1 nfet_05v0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=69745 $Y=46970 $D=2
M10 1 374 ry[7] 1 nfet_05v0 L=6e-07 W=2.724e-05 AD=8.7168e-12 AS=8.7168e-12 PD=3.824e-05 PS=3.824e-05 NRD=0.105727 NRS=0.105727 m=1 nf=3 $X=88785 $Y=46970 $D=2
M11 367 358 2 2 pfet_05v0 L=6e-07 W=2e-05 AD=8.8e-12 AS=8.8e-12 PD=4.088e-05 PS=4.088e-05 NRD=0.022 NRS=0.022 m=1 nf=1 $X=2545 $Y=60125 $D=8
M12 2 371 ly[3] 2 pfet_05v0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=21585 $Y=60125 $D=8
M13 368 361 2 2 pfet_05v0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=24945 $Y=60125 $D=8
M14 365 men 2 2 pfet_05v0 L=6e-07 W=2.275e-06 AD=5.915e-13 AS=1.35362e-12 PD=2.795e-06 PS=5.74e-06 NRD=0.114286 NRS=0.261538 m=1 nf=1 $X=36375 $Y=1335 $D=8
M15 189 clk 365 2 pfet_05v0 L=6e-07 W=2.275e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=37495 $Y=1335 $D=8
M16 366 clk 189 2 pfet_05v0 L=6e-07 W=2.275e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=38615 $Y=1335 $D=8
M17 2 men 366 2 pfet_05v0 L=6e-07 W=2.275e-06 AD=1.34225e-12 AS=5.915e-13 PD=5.73e-06 PS=2.795e-06 NRD=0.259341 NRS=0.114286 m=1 nf=1 $X=39735 $Y=1335 $D=8
M18 2 372 ly[7] 2 pfet_05v0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=43985 $Y=60125 $D=8
M19 369 358 2 2 pfet_05v0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=47345 $Y=60125 $D=8
M20 2 373 ry[3] 2 pfet_05v0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=66385 $Y=60125 $D=8
M21 370 361 2 2 pfet_05v0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=69745 $Y=60125 $D=8
M22 2 374 ry[7] 2 pfet_05v0 L=6e-07 W=6e-05 AD=1.92e-11 AS=1.92e-11 PD=8.192e-05 PS=8.192e-05 NRD=0.048 NRS=0.048 m=1 nf=3 $X=88785 $Y=60125 $D=8
X26 2 188 189 pmos_1p2$$47109164 $T=32795 1405 1 180 $X=28795 $Y=720
X27 1 2 ly[0] 357 ly[1] 359 ly[2] 360 367 371 ICV_21 $T=1275 45270 0 0 $X=1270 $Y=45265
X28 1 2 ly[4] 362 ly[5] 363 ly[6] 364 368 372 ICV_21 $T=23675 45270 0 0 $X=23670 $Y=45265
X29 1 2 ry[0] 357 ry[1] 359 ry[2] 360 369 373 ICV_21 $T=46075 45270 0 0 $X=46070 $Y=45265
X30 1 2 ry[4] 362 ry[5] 363 ry[6] 364 370 374 ICV_21 $T=68475 45270 0 0 $X=68470 $Y=45265
X31 1 195 194 2 192 190 363 364 ICV_22 $T=33645 42985 1 180 $X=28115 $Y=7365
X32 1 195 194 2 193 190 361 362 ICV_22 $T=41810 42985 1 180 $X=36280 $Y=7365
X33 1 195 194 2 192 191 359 360 ICV_22 $T=49980 42985 1 180 $X=44450 $Y=7365
X34 1 195 194 2 193 191 358 357 ICV_22 $T=58150 42985 1 180 $X=52620 $Y=7365
X35 1 190 191 2 A[2] 189 188 ypredec1_bot $T=1920 5135 0 0 $X=1820 $Y=1970
X36 1 192 193 2 A[1] 189 188 ypredec1_bot $T=10375 5135 0 0 $X=10275 $Y=1970
X37 1 194 195 2 A[0] 189 188 ypredec1_bot $T=18830 5135 0 0 $X=18730 $Y=1970
.ENDS
