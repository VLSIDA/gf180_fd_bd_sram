* Subcircuit definition of cell ICV_31
.SUBCKT ICV_31 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49
** N=53 EP=40 IP=82 FDC=220
*.SEEDPROM
M0 7 51 50 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=17060 $D=8
M1 7 53 52 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=18340 $D=8
M2 51 50 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=17060 $D=8
M3 53 52 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=18340 $D=8
X4 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 30 31
+ 32 33 34 35 36 37 38 39 40 41 42 43 44 45
+ ICV_14 $T=-3000 0 1 180 $X=-15340 $Y=-340
X7 7 8 25 26 46 47 50 51 ICV_30 $T=0 0 0 0 $X=-340 $Y=-340
X8 7 8 25 26 52 53 48 49 ICV_30 $T=0 18000 0 0 $X=-340 $Y=17660
.ENDS
