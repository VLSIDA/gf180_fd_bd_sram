* Subcircuit definition of cell xpredec1_bot
.SUBCKT xpredec1_bot 1 2 3 10 11 12 13
** N=32 EP=7 IP=19 FDC=12
X0 1 32 11 10 13 12 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
X2 10 2 32 pmos_1p2$$47337516 $T=3910 18340 0 0 $X=2480 $Y=17635
X3 10 3 2 pmos_1p2$$47337516 $T=6480 18340 0 0 $X=5050 $Y=17635
X4 1 2 32 nmos_1p2$$47336492 $T=3910 36070 0 0 $X=2765 $Y=35385
X5 1 3 2 nmos_1p2$$47336492 $T=6480 36070 0 0 $X=5335 $Y=35385
.ENDS
