* Subcircuit definition of cell wen_wm1
.SUBCKT wen_wm1 vss wep 3 4 5 6 7 8 9 10 11 12 13 men vdd wen GWEN 18 19
** N=43 EP=19 IP=113 FDC=31
M0 3 wen vss vss nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=1765 $Y=5060 $D=2
M1 6 men vss vss nfet_05v0 L=6e-07 W=1.37e-06 AD=3.562e-13 AS=6.028e-13 PD=1.89e-06 PS=3.62e-06 NRD=0.189781 NRS=0.321168 m=1 nf=1 $X=1765 $Y=8905 $D=2
M2 vss GWEN 3 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=2885 $Y=5060 $D=2
M3 vss vss 6 vss nfet_05v0 L=6e-07 W=1.37e-06 AD=6.028e-13 AS=3.562e-13 PD=3.62e-06 PS=1.89e-06 NRD=0.321168 NRS=0.189781 m=1 nf=1 $X=2885 $Y=8905 $D=2
M4 4 3 vss vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=5125 $Y=4650 $D=2
M5 5 6 vss vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=5125 $Y=9315 $D=2
M6 9 6 4 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=7660 $Y=8385 $D=2
M7 7 10 vss vss nfet_05v0 L=6e-07 W=1.37e-06 AD=6.028e-13 AS=6.028e-13 PD=3.62e-06 PS=3.62e-06 NRD=0.321168 NRS=0.321168 m=1 nf=1 $X=8920 $Y=4240 $D=2
M8 11 5 9 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=9970 $Y=9700 $D=2
M9 vss 12 11 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=11090 $Y=9700 $D=2
M10 vss 9 12 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=13330 $Y=9700 $D=2
M11 13 12 vss vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=14450 $Y=9700 $D=2
M12 wep 7 vss vss nfet_05v0 L=6e-07 W=2.4e-06 AD=7.68e-13 AS=7.68e-13 PD=5.12e-06 PS=5.12e-06 NRD=1.2 NRS=1.2 m=1 nf=3 $X=12720 $Y=4810 $D=2
M13 vss 13 8 vss nfet_05v0 L=6e-07 W=1.37e-06 AD=6.028e-13 AS=6.028e-13 PD=3.62e-06 PS=3.62e-06 NRD=0.321168 NRS=0.321168 m=1 nf=1 $X=17810 $Y=9290 $D=2
M14 men 8 10 vss nfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.589e-12 PD=5.58e-06 PS=8.21e-06 NRD=0.229075 NRS=0.30837 m=1 nf=2 $X=20050 $Y=8385 $D=2
M15 vss 13 10 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=22290 $Y=8385 $D=2
M16 18 wen vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=1765 $Y=600 $D=8
M17 19 men vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=1765 $Y=12055 $D=8
M18 3 GWEN 18 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=2885 $Y=600 $D=8
M19 6 vss 19 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=2885 $Y=12055 $D=8
M20 4 3 vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=5125 $Y=600 $D=8
M21 5 6 vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=5125 $Y=12055 $D=8
M22 9 5 4 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=1.17084e-12 AS=9.988e-13 PD=4.78598e-06 PS=5.42e-06 NRD=0.22722 NRS=0.193833 m=1 nf=1 $X=7660 $Y=12055 $D=8
M23 11 6 9 vdd pfet_05v0 L=6e-07 W=9.6e-07 AD=-6.87097e-13 AS=-6.48697e-13 PD=-2.78573e-06 PS=-2.70573e-06 NRD=-0.745548 NRS=-0.703882 m=1 nf=1 $X=9395 $Y=12055 $D=8
M24 vdd 12 11 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=1.14386e-12 PD=5.42e-06 PS=4.72975e-06 NRD=0.193833 NRS=0.221983 m=1 nf=1 $X=11090 $Y=12055 $D=8
M25 vdd 9 12 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=13330 $Y=12055 $D=8
M26 13 12 vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=14450 $Y=12055 $D=8
M27 wep 7 vdd vdd pfet_05v0 L=6e-07 W=6e-06 AD=1.92e-12 AS=1.92e-12 PD=9.92e-06 PS=9.92e-06 NRD=0.48 NRS=0.48 m=1 nf=3 $X=12720 $Y=870 $D=8
M28 men 13 10 vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=20050 $Y=12055 $D=8
X48 vdd 7 10 pfet_05v0_I18 $T=8920 2870 1 0 $X=7880 $Y=540
X49 vdd 8 13 pfet_05v0_I18 $T=16690 12625 0 0 $X=15650 $Y=12005
.ENDS
************* SUBCKT CALLS DEFINITION ***************
.SUBCKT pfet_05v0_I18 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=3.42e-06 AD=8.892e-13 AS=1.5048e-12 PD=4.46e-06 PS=8.6e-06 NRD=0.304094 NRS=0.51462 m=1 nf=2 $X=0 $Y=0 $D=8
.ENDS
