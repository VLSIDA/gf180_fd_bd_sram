* Subcircuit definition of cell gf180mcu_fd_ip_sram__sram64x8m8wm1
.SUBCKT gf180mcu_fd_ip_sram__sram64x8m8wm1 A[5] A[4] A[3] A[2] A[1] A[0] CEN CLK
+ D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] GWEN Q[7] Q[6] Q[5] Q[4] Q[3] Q[2]
+ Q[1] Q[0] VDD VSS WEN[7] WEN[6] WEN[5] WEN[4] WEN[3] WEN[2] WEN[1] WEN[0]
** N=5630 EP=35 IP=395 FDC=6349
M0 VSS 395 599 VSS nfet_05v0 L=6e-07 W=1.36e-06 AD=3.536e-13 AS=5.984e-13 PD=1.88e-06 PS=3.6e-06 NRD=0.191176 NRS=0.323529 m=1 nf=1 $X=233770 $Y=54135 $D=2
M1 599 CLK VSS VSS nfet_05v0 L=6e-07 W=1.36e-06 AD=5.984e-13 AS=3.536e-13 PD=3.6e-06 PS=1.88e-06 NRD=0.323529 NRS=0.191176 m=1 nf=1 $X=234890 $Y=54135 $D=2
M2 592 595 VSS VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=242235 $Y=54135 $D=2
M3 273 598 VSS VSS nfet_05v0 L=1e-06 W=6e-07 AD=2.64e-13 AS=2.64e-13 PD=2.08e-06 PS=2.08e-06 NRD=0.733333 NRS=0.733333 m=1 nf=1 $X=243265 $Y=46010 $D=2
M4 CEN 599 595 VSS nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=245925 $Y=54135 $D=2
M5 242 461 VSS VSS nfet_05v0 L=6e-07 W=4.99e-05 AD=1.47704e-11 AS=1.47704e-11 PD=6.284e-05 PS=6.284e-05 NRD=0.148297 NRS=0.148297 m=1 nf=5 $X=241995 $Y=72320 $D=2
M6 309 273 VSS VSS nfet_05v0 L=6e-07 W=7.5e-07 AD=3.3e-13 AS=3.3e-13 PD=2.38e-06 PS=2.38e-06 NRD=0.586667 NRS=0.586667 m=1 nf=1 $X=246495 $Y=46075 $D=2
M7 346 309 VSS VSS nfet_05v0 L=6e-07 W=3.02e-06 AD=1.3288e-12 AS=1.3288e-12 PD=6.92e-06 PS=6.92e-06 NRD=0.145695 NRS=0.145695 m=1 nf=1 $X=249065 $Y=46070 $D=2
M8 5512 346 VSS VSS nfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=1.34946e-11 PD=2.32e-05 PS=4.655e-05 NRD=0.0114638 NRS=0.0262346 m=1 nf=1 $X=256125 $Y=28435 $D=2
M9 5513 CLK 5512 VSS nfet_05v0 L=6e-07 W=2.268e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=257245 $Y=28435 $D=2
M10 438 592 5513 VSS nfet_05v0 L=6e-07 W=2.268e-05 AD=1.33812e-11 AS=5.8968e-12 PD=4.654e-05 PS=2.32e-05 NRD=0.0260141 NRS=0.0114638 m=1 nf=1 $X=258365 $Y=28435 $D=2
M11 5514 488 VSS VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=4.7177e-12 AS=1.07963e-11 PD=1.8665e-05 PS=3.748e-05 NRD=0.014329 NRS=0.0327914 m=1 nf=1 $X=262120 $Y=29545 $D=2
M12 461 438 5514 VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=263240 $Y=29545 $D=2
M13 5515 438 461 VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=264360 $Y=29545 $D=2
M14 VSS 488 5515 VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=1.07055e-11 AS=4.7177e-12 PD=3.747e-05 PS=1.8665e-05 NRD=0.0325158 NRS=0.014329 m=1 nf=1 $X=265480 $Y=29545 $D=2
M15 5516 461 VSS VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=1.16905e-12 AS=2.7013e-12 PD=5.055e-06 PS=1.027e-05 NRD=0.0567181 NRS=0.131057 m=1 nf=1 $X=268545 $Y=43150 $D=2
M16 488 608 5516 VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=2.27e-14 AS=-2.27e-14 PD=1e-08 PS=-1e-08 NRD=0.00110132 NRS=-0.00110132 m=1 nf=1 $X=269660 $Y=43150 $D=2
M17 5517 608 488 VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=-2.27e-14 AS=2.27e-14 PD=-1e-08 PS=1e-08 NRD=-0.00110132 NRS=0.00110132 m=1 nf=1 $X=270785 $Y=43150 $D=2
M18 VSS 461 5517 VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=2.7013e-12 AS=1.16905e-12 PD=1.027e-05 PS=5.055e-06 NRD=0.131057 NRS=0.0567181 m=1 nf=1 $X=271900 $Y=43150 $D=2
M19 395 242 VSS VSS nfet_05v0 L=6e-07 W=0.0001474 AD=3.8324e-11 AS=4.09772e-11 PD=0.0001578 PS=0.00017326 NRD=0.705563 NRS=0.75441 m=1 nf=20 $X=253180 $Y=76320 $D=2
M20 5594 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=13620 $Y=160970 $D=8
M21 5593 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=13620 $Y=164845 $D=8
M22 5591 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=16720 $Y=160970 $D=8
M23 5592 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=16720 $Y=164845 $D=8
M24 5590 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=19815 $Y=160970 $D=8
M25 5589 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=19815 $Y=164845 $D=8
M26 5587 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=22915 $Y=160970 $D=8
M27 5588 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=22915 $Y=164845 $D=8
M28 5578 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=26005 $Y=160970 $D=8
M29 5577 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=26005 $Y=164845 $D=8
M30 5575 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=29105 $Y=160970 $D=8
M31 5576 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=29105 $Y=164845 $D=8
M32 5580 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=32200 $Y=160970 $D=8
M33 5579 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=32200 $Y=164845 $D=8
M34 625 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=35120 $Y=160970 $D=8
M35 626 5431 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=35120 $Y=164845 $D=8
M36 627 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=38575 $Y=160970 $D=8
M37 628 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=38575 $Y=164845 $D=8
M38 5599 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=41500 $Y=160970 $D=8
M39 5600 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=41500 $Y=164845 $D=8
M40 5598 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=44595 $Y=160970 $D=8
M41 5597 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=44595 $Y=164845 $D=8
M42 5595 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=47695 $Y=160970 $D=8
M43 5596 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=47695 $Y=164845 $D=8
M44 5608 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=50785 $Y=160970 $D=8
M45 5607 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=50785 $Y=164845 $D=8
M46 5605 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=53885 $Y=160970 $D=8
M47 5606 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=53885 $Y=164845 $D=8
M48 5604 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=56980 $Y=160970 $D=8
M49 5603 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=56980 $Y=164845 $D=8
M50 5601 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=60080 $Y=160970 $D=8
M51 5602 5432 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=60080 $Y=164845 $D=8
M52 5616 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=67620 $Y=160970 $D=8
M53 5615 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=67620 $Y=164845 $D=8
M54 5613 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=70720 $Y=160970 $D=8
M55 5614 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=70720 $Y=164845 $D=8
M56 5612 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=73815 $Y=160970 $D=8
M57 5611 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=73815 $Y=164845 $D=8
M58 5609 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=76915 $Y=160970 $D=8
M59 5610 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=76915 $Y=164845 $D=8
M60 5584 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=80005 $Y=160970 $D=8
M61 5583 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=80005 $Y=164845 $D=8
M62 5581 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=83105 $Y=160970 $D=8
M63 5582 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=83105 $Y=164845 $D=8
M64 5586 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=86200 $Y=160970 $D=8
M65 5585 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=86200 $Y=164845 $D=8
M66 629 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=89120 $Y=160970 $D=8
M67 630 5433 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=89120 $Y=164845 $D=8
M68 631 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=92575 $Y=160970 $D=8
M69 632 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=92575 $Y=164845 $D=8
M70 5629 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=95500 $Y=160970 $D=8
M71 5630 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=95500 $Y=164845 $D=8
M72 5628 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=98595 $Y=160970 $D=8
M73 5627 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=98595 $Y=164845 $D=8
M74 5625 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=101695 $Y=160970 $D=8
M75 5626 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=101695 $Y=164845 $D=8
M76 5624 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=104785 $Y=160970 $D=8
M77 5623 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=104785 $Y=164845 $D=8
M78 5621 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=107885 $Y=160970 $D=8
M79 5622 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=107885 $Y=164845 $D=8
M80 5620 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=110980 $Y=160970 $D=8
M81 5619 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=110980 $Y=164845 $D=8
M82 5617 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=114080 $Y=160970 $D=8
M83 5618 5434 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=114080 $Y=164845 $D=8
M84 5518 395 VDD VDD pfet_05v0 L=5.95e-07 W=2.28e-06 AD=5.985e-13 AS=1.3566e-12 PD=2.805e-06 PS=5.75e-06 NRD=0.115132 NRS=0.260965 m=1 nf=1 $X=233770 $Y=57780 $D=8
M85 593 599 VDD VDD pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=233770 $Y=63100 $D=8
M86 599 CLK 5518 VDD pfet_05v0 L=5.95e-07 W=2.28e-06 AD=1.3566e-12 AS=5.985e-13 PD=5.75e-06 PS=2.805e-06 NRD=0.260965 NRS=0.115132 m=1 nf=1 $X=234890 $Y=57780 $D=8
M87 592 595 VDD VDD pfet_05v0 L=6e-07 W=1.134e-05 AD=2.9484e-12 AS=4.9896e-12 PD=1.238e-05 PS=2.444e-05 NRD=0.0917108 NRS=0.155203 m=1 nf=2 $X=242235 $Y=57810 $D=8
M88 273 598 VDD VDD pfet_05v0 L=1e-06 W=9e-07 AD=3.96e-13 AS=3.96e-13 PD=2.68e-06 PS=2.68e-06 NRD=0.488889 NRS=0.488889 m=1 nf=1 $X=243265 $Y=42525 $D=8
M89 CEN 593 595 VDD pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=245925 $Y=59010 $D=8
M90 594 599 595 VDD pfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=245925 $Y=64875 $D=8
M91 309 273 VDD VDD pfet_05v0 L=6e-07 W=1.89e-06 AD=8.316e-13 AS=8.316e-13 PD=4.66e-06 PS=4.66e-06 NRD=0.232804 NRS=0.232804 m=1 nf=1 $X=246495 $Y=41535 $D=8
M92 346 309 VDD VDD pfet_05v0 L=6e-07 W=7.54e-06 AD=1.9604e-12 AS=3.3176e-12 PD=8.58e-06 PS=1.684e-05 NRD=0.137931 NRS=0.233422 m=1 nf=2 $X=249065 $Y=39655 $D=8
M93 242 461 VDD VDD pfet_05v0 L=6e-07 W=0.0001248 AD=3.2448e-11 AS=3.69283e-11 PD=0.00013 PS=0.000130718 NRD=0.208333 NRS=0.237099 m=1 nf=10 $X=240535 $Y=94430 $D=8
M94 438 346 VDD VDD pfet_05v0 L=6e-07 W=1.95e-05 AD=5.07e-12 AS=8.58e-12 PD=2.002e-05 PS=3.988e-05 NRD=0.0133333 NRS=0.0225641 m=1 nf=1 $X=256125 $Y=53590 $D=8
M95 VDD CLK 438 VDD pfet_05v0 L=6e-07 W=1.95e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=257245 $Y=53590 $D=8
M96 438 592 VDD VDD pfet_05v0 L=6e-07 W=1.95e-05 AD=8.58e-12 AS=5.07e-12 PD=3.988e-05 PS=2.002e-05 NRD=0.0225641 NRS=0.0133333 m=1 nf=1 $X=258365 $Y=53590 $D=8
M97 VDD 488 461 VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=9.9792e-12 PD=2.32e-05 PS=4.624e-05 NRD=0.0114638 NRS=0.0194004 m=1 nf=1 $X=262120 $Y=50420 $D=8
M98 461 438 VDD VDD pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.64e-05 PS=4.64e-05 NRD=0.0229277 NRS=0.0229277 m=1 nf=2 $X=263240 $Y=50420 $D=8
M99 461 488 VDD VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=9.9792e-12 AS=5.8968e-12 PD=4.624e-05 PS=2.32e-05 NRD=0.0194004 NRS=0.0114638 m=1 nf=1 $X=265480 $Y=50420 $D=8
M100 VDD 461 488 VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=9.9792e-12 PD=2.32e-05 PS=4.624e-05 NRD=0.0114638 NRS=0.0194004 m=1 nf=1 $X=268545 $Y=50420 $D=8
M101 488 608 VDD VDD pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.64e-05 PS=4.64e-05 NRD=0.0229277 NRS=0.0229277 m=1 nf=2 $X=269665 $Y=50420 $D=8
M102 488 461 VDD VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=9.9792e-12 AS=5.8968e-12 PD=4.624e-05 PS=2.32e-05 NRD=0.0194004 NRS=0.0114638 m=1 nf=1 $X=271905 $Y=50420 $D=8
M103 395 242 VDD VDD pfet_05v0 L=6e-07 W=0.0003674 AD=9.5524e-11 AS=1.02119e-10 PD=0.0003778 PS=0.000378518 NRD=0.28307 NRS=0.302613 m=1 nf=20 $X=253180 $Y=88540 $D=8
M104 5566 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=311500 $Y=160970 $D=8
M105 5565 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=311500 $Y=164845 $D=8
M106 5563 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=314600 $Y=160970 $D=8
M107 5564 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=314600 $Y=164845 $D=8
M108 5562 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=317695 $Y=160970 $D=8
M109 5561 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=317695 $Y=164845 $D=8
M110 5559 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=320795 $Y=160970 $D=8
M111 5560 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=320795 $Y=164845 $D=8
M112 5550 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=323885 $Y=160970 $D=8
M113 5549 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=323885 $Y=164845 $D=8
M114 5547 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=326985 $Y=160970 $D=8
M115 5548 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=326985 $Y=164845 $D=8
M116 5552 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=330080 $Y=160970 $D=8
M117 5551 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=330080 $Y=164845 $D=8
M118 617 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=333000 $Y=160970 $D=8
M119 618 5428 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=333000 $Y=164845 $D=8
M120 619 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=336455 $Y=160970 $D=8
M121 620 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=336455 $Y=164845 $D=8
M122 5523 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=339380 $Y=160970 $D=8
M123 5524 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=339380 $Y=164845 $D=8
M124 5522 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=342475 $Y=160970 $D=8
M125 5521 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=342475 $Y=164845 $D=8
M126 5519 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=345575 $Y=160970 $D=8
M127 5520 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=345575 $Y=164845 $D=8
M128 5532 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=348665 $Y=160970 $D=8
M129 5531 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=348665 $Y=164845 $D=8
M130 5529 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=351765 $Y=160970 $D=8
M131 5530 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=351765 $Y=164845 $D=8
M132 5528 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=354860 $Y=160970 $D=8
M133 5527 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=354860 $Y=164845 $D=8
M134 5525 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=357960 $Y=160970 $D=8
M135 5526 5429 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=357960 $Y=164845 $D=8
M136 5574 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=365500 $Y=160970 $D=8
M137 5573 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=365500 $Y=164845 $D=8
M138 5571 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=368600 $Y=160970 $D=8
M139 5572 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=368600 $Y=164845 $D=8
M140 5570 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=371695 $Y=160970 $D=8
M141 5569 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=371695 $Y=164845 $D=8
M142 5567 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=374795 $Y=160970 $D=8
M143 5568 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=374795 $Y=164845 $D=8
M144 5556 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=377885 $Y=160970 $D=8
M145 5555 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=377885 $Y=164845 $D=8
M146 5553 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=380985 $Y=160970 $D=8
M147 5554 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=380985 $Y=164845 $D=8
M148 5558 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=384080 $Y=160970 $D=8
M149 5557 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=384080 $Y=164845 $D=8
M150 621 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=387000 $Y=160970 $D=8
M151 622 5430 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=387000 $Y=164845 $D=8
M152 623 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=390455 $Y=160970 $D=8
M153 624 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=390455 $Y=164845 $D=8
M154 5537 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=393380 $Y=160970 $D=8
M155 5538 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=393380 $Y=164845 $D=8
M156 5536 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=396475 $Y=160970 $D=8
M157 5535 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=396475 $Y=164845 $D=8
M158 5533 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=399575 $Y=160970 $D=8
M159 5534 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=399575 $Y=164845 $D=8
M160 5546 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=402665 $Y=160970 $D=8
M161 5545 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=402665 $Y=164845 $D=8
M162 5543 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=405765 $Y=160970 $D=8
M163 5544 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=405765 $Y=164845 $D=8
M164 5542 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=408860 $Y=160970 $D=8
M165 5541 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=408860 $Y=164845 $D=8
M166 5539 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=411960 $Y=160970 $D=8
M167 5540 616 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=411960 $Y=164845 $D=8
X175 VSS 593 599 VSS nmos_1p2$$46563372 $T=233925 66830 0 0 $X=232780 $Y=66145
X176 594 VSS 592 VSS nmos_1p2$$46563372 $T=243510 68190 1 0 $X=242365 $Y=66555
X177 595 594 593 VSS nmos_1p2$$46563372 $T=246080 68190 1 0 $X=244935 $Y=66555
X178 VDD 594 592 pmos_1p2$$46273580 $T=242390 65835 1 0 $X=240960 $Y=64015
X180 VSS 608 616 VDD 5452 WEN[5] 5429 619 620 395 WEN[7] 623 624 WEN[4] 5428 617 618 WEN[6] 5430 621
+ 622 5461 5462 5463 5464 5465 5466 5467 5468 607 5451 5459 5460 5458 5457 5456 5455 5454 5453 D[5]
+ Q[5] D[7] Q[7] D[4] Q[4] D[6] Q[6] 5519 5520 5521 5522 5523 5524 5525 5526 5527 5528 5529 5530 5531
+ 5532 5533 5534 5535 5536 5537 5538 5539 5540 5541 5542 5543 5544 5545 5546 5547 5548 5549 5550 5551
+ 5552 5553 5554 5555 5556 5557 5558 5559 5560 5561 5562 5563 5564 5565 5566 5567 5568 5569 5570 5571
+ 5572 5573 5574
+ rcol4_64 $T=302555 25095 0 0 $X=297105 $Y=5955
X191 VSS 597 CLK nfet_05v0_I09 $T=234280 46585 1 0 $X=233600 $Y=45365
X192 VSS 598 597 nfet_05v0_I09 $T=239670 46585 1 0 $X=238990 $Y=45365
X193 VDD 597 CLK pfet_05v0_I15 $T=234280 43425 1 0 $X=233240 $Y=41905
X194 VDD 598 597 pfet_05v0_I15 $T=239670 43425 1 0 $X=238630 $Y=41905
X197 VSS 395 VDD CLK A[5] A[4] A[3] 5496 5497 5498 5499 5500 5501 5502 5503 xpredec1 $T=219860 111460 0 0 $X=219855 $Y=111455
X198 VSS 5450 VDD GWEN CLK 5451 607 wen_v2 $T=208415 16605 0 0 $X=208280 $Y=15275
X201 VSS VDD 395 CLK VSS VSS 5485 5486 5490 5491 xpredec0 $T=146075 111460 0 0 $X=144630 $Y=111455
X202 VSS VDD 395 CLK VSS VSS 5492 5493 5494 5495 xpredec0 $T=182970 111460 0 0 $X=181525 $Y=111455
X203 VSS VDD 395 CLK 5448 5449 5442 5443 5444 5445 5446 5447 5460 5459 5458 5457 5456 5455 5454 5453
+ A[2] A[1] A[0]
+ ypredec1 $T=145470 26355 0 0 $X=146365 $Y=26735
X205 395 VSS 5452 VDD 5503 5502 5501 5500 5499 5498 5497 5496 5469 5470 5471 5472 5473 5474 5475 5476
+ 5462 5463 5465 5467 5468 5464 5466 5461
+ xdec8_64 $T=143385 180635 0 0 $X=126565 $Y=178920
X206 VSS VDD WEN[1] 5432 627 628 395 WEN[3] 5434 631 632 WEN[0] 5431 625 626 WEN[2] 5433 629 630 5469
+ 5470 5471 5472 5473 5474 5475 5476 5451 607 5442 5443 5444 5445 5446 5447 5448 5449 D[1] Q[1] D[3]
+ Q[3] D[0] Q[0] D[2] Q[2] 5575 5576 5577 5578 5579 5580 5581 5582 5583 5584 5585 5586 5587 5588 5589
+ 5590 5591 5592 5593 5594 5595 5596 5597 5598 5599 5600 5601 5602 5603 5604 5605 5606 5607 5608 5609
+ 5610 5611 5612 5613 5614 5615 5616 5617 5618 5619 5620 5621 5622 5623 5624 5625 5626 5627 5628 5629
+ 5630
+ lcol4_64 $T=14605 25095 0 0 $X=2855 $Y=4030
.ENDS
