* Subcircuit definition of cell 018SRAM_cell1_dummy_R
.SUBCKT 018SRAM_cell1_dummy_R
** N=8 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
