* Subcircuit definition of cell nmos_1p2$$46551084
.SUBCKT nmos_1p2$$46551084
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
