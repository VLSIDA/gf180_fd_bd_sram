* Subcircuit definition of cell nmos_1p2$$47342636
.SUBCKT nmos_1p2$$47342636
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
