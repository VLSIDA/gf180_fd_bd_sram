* Subcircuit definition of cell xdec8_64
.SUBCKT xdec8_64 men vss DRWL vdd xa[0] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] xa[7] LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] LWL[6] LWL[7]
+ RWL[1] RWL[2] RWL[4] RWL[6] RWL[7] RWL[3] RWL[5] RWL[0]
** N=317 EP=28 IP=541 FDC=156
M0 vss 288 LWL[0] vss nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=24970 $Y=260 $D=2
M1 288 272 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=24970 $Y=2660 $D=2
M2 vss 270 286 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=24970 $Y=5740 $D=2
M3 vss 286 LWL[1] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=24970 $Y=7020 $D=2
M4 vss 292 LWL[2] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=24970 $Y=9260 $D=2
M5 292 276 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=24970 $Y=11660 $D=2
M6 vss 274 290 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=24970 $Y=14740 $D=2
M7 vss 290 LWL[3] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=24970 $Y=16020 $D=2
M8 vss 296 LWL[4] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=24970 $Y=18260 $D=2
M9 296 280 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=24970 $Y=20660 $D=2
M10 vss 278 294 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=24970 $Y=23740 $D=2
M11 vss 294 LWL[5] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=24970 $Y=25020 $D=2
M12 vss 300 LWL[6] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=24970 $Y=27260 $D=2
M13 300 284 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=24970 $Y=29660 $D=2
M14 vss 282 298 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=24970 $Y=32740 $D=2
M15 vss 298 LWL[7] vss nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=24970 $Y=34020 $D=2
M16 272 273 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=55250 $Y=260 $D=2
M17 vss 271 270 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=55250 $Y=8140 $D=2
M18 276 277 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=55250 $Y=9260 $D=2
M19 vss 275 274 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=55250 $Y=17140 $D=2
M20 280 281 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=55250 $Y=18260 $D=2
M21 vss 279 278 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=55250 $Y=26140 $D=2
M22 284 285 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=55250 $Y=27260 $D=2
M23 vss 283 282 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=55250 $Y=35140 $D=2
M24 29 vdd men vss nfet_05v0 L=6e-07 W=6.59e-06 AD=2.8996e-12 AS=2.8996e-12 PD=1.406e-05 PS=1.406e-05 NRD=0.0667678 NRS=0.0667678 m=1 nf=1 $X=61430 $Y=38365 $D=2
M25 305 vdd vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=7.32375e-13 AS=2.079e-12 PD=3.615e-06 PS=7.62e-06 NRD=0.0738095 NRS=0.209524 m=1 nf=1 $X=75090 $Y=315 $D=2
M26 304 vdd 305 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=75090 $Y=1380 $D=2
M27 273 xa[0] 304 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=75090 $Y=2500 $D=2
M28 302 xa[1] 271 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=75090 $Y=5900 $D=2
M29 303 vdd 302 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=75090 $Y=7020 $D=2
M30 vss vdd 303 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=75090 $Y=8085 $D=2
M31 309 vdd vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=75090 $Y=9315 $D=2
M32 308 vdd 309 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=75090 $Y=10380 $D=2
M33 277 xa[2] 308 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=75090 $Y=11500 $D=2
M34 306 xa[3] 275 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=75090 $Y=14900 $D=2
M35 307 vdd 306 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=75090 $Y=16020 $D=2
M36 vss vdd 307 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=75090 $Y=17085 $D=2
M37 313 vdd vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=75090 $Y=18315 $D=2
M38 312 vdd 313 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=75090 $Y=19380 $D=2
M39 281 xa[4] 312 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=75090 $Y=20500 $D=2
M40 310 xa[5] 279 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=75090 $Y=23900 $D=2
M41 311 vdd 310 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=75090 $Y=25020 $D=2
M42 vss vdd 311 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=75090 $Y=26085 $D=2
M43 317 vdd vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=75090 $Y=27315 $D=2
M44 316 vdd 317 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=75090 $Y=28380 $D=2
M45 285 xa[6] 316 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=75090 $Y=29500 $D=2
M46 314 xa[7] 283 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=75090 $Y=32900 $D=2
M47 315 vdd 314 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=75090 $Y=34020 $D=2
M48 vss vdd 315 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.079e-12 AS=7.32375e-13 PD=7.62e-06 PS=3.615e-06 NRD=0.209524 NRS=0.0738095 m=1 nf=1 $X=75090 $Y=35085 $D=2
M49 vss 289 RWL[0] vss nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=108885 $Y=260 $D=2
M50 289 272 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=108885 $Y=2660 $D=2
M51 vss 270 287 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=108885 $Y=5740 $D=2
M52 vss 287 RWL[1] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=108885 $Y=7020 $D=2
M53 vss 293 RWL[2] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=108885 $Y=9260 $D=2
M54 293 276 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=108885 $Y=11660 $D=2
M55 vss 274 291 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=108885 $Y=14740 $D=2
M56 vss 291 RWL[3] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=108885 $Y=16020 $D=2
M57 vss 297 RWL[4] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=108885 $Y=18260 $D=2
M58 297 280 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=108885 $Y=20660 $D=2
M59 vss 278 295 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=108885 $Y=23740 $D=2
M60 vss 295 RWL[5] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=108885 $Y=25020 $D=2
M61 vss 301 RWL[6] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=108885 $Y=27260 $D=2
M62 301 284 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=108885 $Y=29660 $D=2
M63 vss 282 299 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=108885 $Y=32740 $D=2
M64 vss 299 RWL[7] vss nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=108885 $Y=34020 $D=2
M65 vdd vss vdd vdd pfet_05v0 L=3.94e-06 W=4.9455e-05 AD=0 AS=3.14863e-11 PD=0 PS=0.00012136 NRD=0 NRS=1.04277 m=1 nf=9 $X=2985 $Y=280 $D=8
M66 vdd 288 LWL[0] vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=13295 $Y=260 $D=8
M67 LWL[1] 286 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=13295 $Y=5900 $D=8
M68 vdd 292 LWL[2] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=13295 $Y=9260 $D=8
M69 LWL[3] 290 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=13295 $Y=14900 $D=8
M70 vdd 296 LWL[4] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=13295 $Y=18260 $D=8
M71 LWL[5] 294 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=13295 $Y=23900 $D=8
M72 vdd 300 LWL[6] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=13295 $Y=27260 $D=8
M73 LWL[7] 298 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=13295 $Y=32900 $D=8
M74 vdd vdd 273 vdd pfet_05v0 L=6e-07 W=5.24e-06 AD=1.834e-12 AS=1.3624e-12 PD=9.26e-06 PS=6.28e-06 NRD=0.267176 NRS=0.198473 m=1 nf=2 $X=80610 $Y=260 $D=8
M75 273 xa[0] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=80610 $Y=2500 $D=8
M76 vdd xa[1] 271 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=80610 $Y=5900 $D=8
M77 vdd vdd 271 vdd pfet_05v0 L=6e-07 W=5.24e-06 AD=1.3624e-12 AS=1.3624e-12 PD=6.28e-06 PS=6.28e-06 NRD=0.198473 NRS=0.198473 m=1 nf=2 $X=80610 $Y=7020 $D=8
M78 vdd vdd 277 vdd pfet_05v0 L=6e-07 W=5.24e-06 AD=1.3624e-12 AS=1.3624e-12 PD=6.28e-06 PS=6.28e-06 NRD=0.198473 NRS=0.198473 m=1 nf=2 $X=80610 $Y=9260 $D=8
M79 277 xa[2] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=80610 $Y=11500 $D=8
M80 vdd xa[3] 275 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=80610 $Y=14900 $D=8
M81 vdd vdd 275 vdd pfet_05v0 L=6e-07 W=5.24e-06 AD=1.3624e-12 AS=1.3624e-12 PD=6.28e-06 PS=6.28e-06 NRD=0.198473 NRS=0.198473 m=1 nf=2 $X=80610 $Y=16020 $D=8
M82 vdd vdd 281 vdd pfet_05v0 L=6e-07 W=5.24e-06 AD=1.3624e-12 AS=1.3624e-12 PD=6.28e-06 PS=6.28e-06 NRD=0.198473 NRS=0.198473 m=1 nf=2 $X=80610 $Y=18260 $D=8
M83 281 xa[4] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=80610 $Y=20500 $D=8
M84 vdd xa[5] 279 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=80610 $Y=23900 $D=8
M85 vdd vdd 279 vdd pfet_05v0 L=6e-07 W=5.24e-06 AD=1.3624e-12 AS=1.3624e-12 PD=6.28e-06 PS=6.28e-06 NRD=0.198473 NRS=0.198473 m=1 nf=2 $X=80610 $Y=25020 $D=8
M86 vdd vdd 285 vdd pfet_05v0 L=6e-07 W=5.24e-06 AD=1.3624e-12 AS=1.3624e-12 PD=6.28e-06 PS=6.28e-06 NRD=0.198473 NRS=0.198473 m=1 nf=2 $X=80610 $Y=27260 $D=8
M87 285 xa[6] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=80610 $Y=29500 $D=8
M88 vdd xa[7] 283 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=80610 $Y=32900 $D=8
M89 vdd vdd 283 vdd pfet_05v0 L=6e-07 W=5.24e-06 AD=1.834e-12 AS=1.3624e-12 PD=9.26e-06 PS=6.28e-06 NRD=0.267176 NRS=0.198473 m=1 nf=2 $X=80610 $Y=34020 $D=8
M90 vdd 289 RWL[0] vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=115560 $Y=260 $D=8
M91 RWL[1] 287 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=115560 $Y=5900 $D=8
M92 vdd 293 RWL[2] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=115560 $Y=9260 $D=8
M93 RWL[3] 291 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=115560 $Y=14900 $D=8
M94 vdd 297 RWL[4] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=115560 $Y=18260 $D=8
M95 RWL[5] 295 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=115560 $Y=23900 $D=8
M96 vdd 301 RWL[6] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=115560 $Y=27260 $D=8
M97 RWL[7] 299 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=115560 $Y=32900 $D=8
M98 vdd vss vdd vdd pfet_05v0 L=3.94e-06 W=4.9455e-05 AD=0 AS=3.14863e-11 PD=0 PS=0.00012136 NRD=0 NRS=1.04277 m=1 nf=9 $X=130365 $Y=280 $D=8
X110 DLWL vss 37 nfet_05v0_I14 $T=31730 38360 0 90 $X=21000 $Y=37680
X111 DRWL vss 38 nfet_05v0_I14 $T=116730 38360 0 90 $X=106000 $Y=37680
X112 vdd DLWL 37 pmos_1p2$$204216364_R90 $T=46225 38515 0 90 $X=32935 $Y=37035
X113 vdd DRWL 38 pmos_1p2$$204216364_R90 $T=104750 38515 0 90 $X=91460 $Y=37035
X114 37 vdd 29 vdd pfet_05v0_I03 $T=55020 38360 0 90 $X=47810 $Y=37320
X115 men 29 vss vdd pfet_05v0_I03 $T=76520 38360 0 90 $X=69310 $Y=37320
X116 38 vdd 29 vdd pfet_05v0_I03 $T=89870 38360 0 90 $X=82660 $Y=37320
X117 37 vss 29 nfet_05v0_I05 $T=59565 38360 0 90 $X=56305 $Y=37680
X118 38 vss 29 nfet_05v0_I05 $T=81415 38360 0 90 $X=78155 $Y=37680
X119 vss vdd 270 men 271 272 273 286 287 288 289 ICV_24 $T=8635 4500 1 0 $X=8630 $Y=-1140
X120 vss vdd 274 men 275 276 277 290 291 292 293 ICV_24 $T=8635 13500 1 0 $X=8630 $Y=7860
X121 vss vdd 278 men 279 280 281 294 295 296 297 ICV_24 $T=8635 22500 1 0 $X=8630 $Y=16860
X122 vss vdd 282 men 283 284 285 298 299 300 301 ICV_24 $T=8635 31500 1 0 $X=8630 $Y=25860
.ENDS
