* Subcircuit definition of cell M1_PSUB_I04
.SUBCKT M1_PSUB_I04
** N=2401 EP=0 IP=0 FDC=0
.ENDS
