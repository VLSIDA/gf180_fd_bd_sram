* Subcircuit definition of cell ICV_10
.SUBCKT ICV_10
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
