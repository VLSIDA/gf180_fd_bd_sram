* Subcircuit definition of cell M1_PSUB_I04
.SUBCKT M1_PSUB_I04
** N=3805 EP=0 IP=0 FDC=0
.ENDS
