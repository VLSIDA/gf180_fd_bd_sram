* Subcircuit definition of cell M1_PSUB_I01
.SUBCKT M1_PSUB_I01
** N=666 EP=0 IP=0 FDC=0
.ENDS
