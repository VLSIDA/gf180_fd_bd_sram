* Subcircuit definition of cell nfet_05v0_I15
.SUBCKT nfet_05v0_I15
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
