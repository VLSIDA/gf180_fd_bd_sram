* Subcircuit definition of cell ypass_gate
.SUBCKT ypass_gate vss 3 b d bb db ypass pcb vdd
** N=26 EP=9 IP=25 FDC=5
*.SEEDPROM
X2 bb b pcb vdd pfet_05v0_I09 $T=1240 50985 1 0 $X=200 $Y=43555
X3 bb db 3 vdd pfet_05v0_I09 $T=1250 43050 1 0 $X=210 $Y=35620
X4 b d 3 vdd pmos_1p2$$46889004 $T=1405 15300 1 0 $X=-25 $Y=7790
X5 b d ypass vss nmos_1p2$$47119404 $T=1405 24575 1 0 $X=260 $Y=17090
X6 bb db ypass vss nmos_1p2$$47119404 $T=1405 34595 1 0 $X=260 $Y=27110
.ENDS
************* SUBCKT CALLS DEFINITION ***************
.SUBCKT pfet_05v0_I09 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 pfet_05v0 L=6e-07 W=6.81e-06 AD=2.9964e-12 AS=2.9964e-12 PD=1.45e-05 PS=1.45e-05 NRD=0.0646109 NRS=0.0646109 m=1 nf=1 $X=0 $Y=0 $D=8
.ENDS
.SUBCKT pmos_1p2$$46889004 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
X0 1 2 3 4 pfet_05v0_I09 $T=-155 0 0 0 $X=-1195 $Y=-620
.ENDS
.SUBCKT nmos_1p2$$47119404 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
X0 1 2 3 4 nfet_05v0_I12 $T=-155 0 0 0 $X=-835 $Y=-620
.ENDS
.SUBCKT nfet_05v0_I12 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nfet_05v0 L=6e-07 W=6.81e-06 AD=2.9964e-12 AS=2.9964e-12 PD=1.45e-05 PS=1.45e-05 NRD=0.0646109 NRS=0.0646109 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
