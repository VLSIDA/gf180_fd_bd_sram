* Subcircuit definition of cell pfet_05v0_I08
.SUBCKT pfet_05v0_I08 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=1.2e-06 W=9e-07 AD=3.96e-13 AS=3.96e-13 PD=2.68e-06 PS=2.68e-06 NRD=0.488889 NRS=0.488889 m=1 nf=1 $X=0 $Y=0 $D=8
.ENDS
