* Subcircuit definition of cell nfet_05v0_I17
.SUBCKT nfet_05v0_I17 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nfet_05v0 L=6e-07 W=1.135e-05 AD=3.3596e-12 AS=3.3596e-12 PD=1.658e-05 PS=1.658e-05 NRD=0.651982 NRS=0.651982 m=1 nf=5 $X=0 $Y=0 $D=2
.ENDS
