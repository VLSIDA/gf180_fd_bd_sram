* Subcircuit definition of cell ICV_29
.SUBCKT ICV_29 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
** N=30 EP=30 IP=36 FDC=80
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 15 16 17 18 19 20 21 22 ICV_28 $T=0 0 0 0 $X=-340 $Y=-340
X1 1 2 3 4 5 6 11 12 13 14 23 24 25 26 27 28 29 30 ICV_28 $T=6000 0 0 0 $X=5660 $Y=-340
.ENDS
