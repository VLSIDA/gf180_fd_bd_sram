* Subcircuit definition of cell ICV_17
.SUBCKT ICV_17 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 33 34 35 36 37 38 39 40
** N=40 EP=34 IP=50 FDC=176
*.SEEDPROM
X0 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ ICV_14 $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
