* Subcircuit definition of cell M1_NWELL_I02
.SUBCKT M1_NWELL_I02
** N=4 EP=0 IP=0 FDC=0
.ENDS
