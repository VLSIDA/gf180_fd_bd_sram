* Subcircuit definition of cell ICV_25
.SUBCKT ICV_25 1 2 7 8 9 10 11 12
** N=16 EP=8 IP=20 FDC=20
*.SEEDPROM
M0 1 14 13 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=-5440 $D=8
M1 1 16 15 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=-4160 $D=8
M2 14 13 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=-5440 $D=8
M3 16 15 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=-4160 $D=8
X4 7 8 2 9 10 13 14 ICV_24 $T=0 -9000 0 0 $X=-340 $Y=-13840
X5 7 8 2 15 16 11 12 ICV_24 $T=0 0 0 0 $X=-340 $Y=-4840
.ENDS
