* Subcircuit definition of cell ICV_10
.SUBCKT ICV_10 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36 37 38
** N=54 EP=34 IP=57 FDC=32
*.SEEDPROM
X0 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 ICV_8 $T=-15000 0 0 0 $X=-24340 $Y=-340
X1 4 6 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 ICV_9 $T=0 0 0 0 $X=-12340 $Y=-340
.ENDS
