* Subcircuit definition of cell xpredec0_bot
.SUBCKT xpredec0_bot 1 2 3 8 9 10 11
** N=33 EP=7 IP=7 FDC=12
M0 2 33 1 1 nfet_05v0 L=6e-07 W=7.04e-06 AD=3.0976e-12 AS=3.0976e-12 PD=1.496e-05 PS=1.496e-05 NRD=0.0625 NRS=0.0625 m=1 nf=1 $X=3755 $Y=35615 $D=2
M1 3 2 1 1 nfet_05v0 L=6e-07 W=5.22e-06 AD=2.2968e-12 AS=2.2968e-12 PD=1.132e-05 PS=1.132e-05 NRD=0.0842912 NRS=0.0842912 m=1 nf=1 $X=6325 $Y=36010 $D=2
M2 2 33 8 8 pfet_05v0 L=6e-07 W=1.769e-05 AD=7.7836e-12 AS=7.7836e-12 PD=3.626e-05 PS=3.626e-05 NRD=0.0248728 NRS=0.0248728 m=1 nf=1 $X=3755 $Y=16320 $D=8
M3 3 2 8 8 pfet_05v0 L=6e-07 W=1.316e-05 AD=5.7904e-12 AS=5.7904e-12 PD=2.72e-05 PS=2.72e-05 NRD=0.0334347 NRS=0.0334347 m=1 nf=1 $X=6325 $Y=20855 $D=8
X4 1 33 9 8 11 10 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
.ENDS
************* SUBCKT CALLS DEFINITION ***************
.SUBCKT alatch vss ab a vdd enb en
** N=16 EP=6 IP=24 FDC=8
M0 ab 12 vss vss nfet_05v0 L=6e-07 W=3.64e-06 AD=9.464e-13 AS=1.6016e-12 PD=4.68e-06 PS=9.04e-06 NRD=0.285714 NRS=0.483516 m=1 nf=2 $X=2590 $Y=1475 $D=2
M1 vss ab 11 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=3710 $Y=12935 $D=2
M2 a en 12 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=6280 $Y=1020 $D=2
M3 11 enb 12 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=6280 $Y=12935 $D=2
M4 ab 12 vdd vdd pfet_05v0 L=6e-07 W=9.08e-06 AD=2.3608e-12 AS=3.9952e-12 PD=1.012e-05 PS=1.992e-05 NRD=0.114537 NRS=0.193833 m=1 nf=2 $X=2590 $Y=4695 $D=8
M5 a enb 12 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=6280 $Y=5895 $D=8
X10 11 vdd ab vdd pmos_1p2$$47330348_161 $T=3865 11540 1 0 $X=2435 $Y=9910
X11 12 11 en vdd pmos_1p2$$47330348_161 $T=6435 11540 1 0 $X=5005 $Y=9910
.ENDS
.SUBCKT pmos_1p2$$47330348_161 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
M0 2 3 1 4 pfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
