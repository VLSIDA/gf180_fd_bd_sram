* Subcircuit definition of cell ICV_18
.SUBCKT ICV_18 7 8 13 14 18 19 20 21
** N=25 EP=8 IP=32 FDC=20
*.SEEDPROM
M0 7 23 22 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=8060 $D=8
M1 7 25 24 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=9340 $D=8
M2 23 22 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=8060 $D=8
M3 25 24 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=9340 $D=8
X4 8 13 14 18 22 19 23 ICV_17 $T=0 0 0 0 $X=-3340 $Y=-340
X5 8 13 14 24 20 25 21 ICV_17 $T=0 9000 0 0 $X=-3340 $Y=8660
.ENDS
