* Subcircuit definition of cell ICV_7
.SUBCKT ICV_7 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 48
+ 80 112 144
** N=175 EP=43 IP=215 FDC=392
*.SEEDPROM
M0 2 111 79 2 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=143060 $D=8
M1 2 43 41 2 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=144340 $D=8
M2 111 79 2 2 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=143060 $D=8
M3 43 41 2 2 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=144340 $D=8
M4 2 175 143 2 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=143060 $D=8
M5 2 47 45 2 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=144340 $D=8
M6 175 143 2 2 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=143060 $D=8
M7 47 45 2 2 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=144340 $D=8
X8 1 3 40 41 42 43 44 45 46 47 ICV_6 $T=0 148500 1 0 $X=-3340 $Y=143660
X9 2 1 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 48 36 49 50 51 52
+ 53 54 55 37 80 81 82 83 84 85 86 87 56 57 58 59 60 61 62 63
+ 88 89 90 91 92 93 94 95 64 65 66 67 68 69 70 71 96 97 98 99
+ 100 101 102 103 72 73 74 75 76 77 78 79 104 105 106 107 108 109 110 111
+ Cell_array32x1 $T=-3000 0 0 0 $X=-3340 $Y=-340
X10 2 1 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 112 38 113 114 115 116
+ 117 118 119 39 144 145 146 147 148 149 150 151 120 121 122 123 124 125 126 127
+ 152 153 154 155 156 157 158 159 128 129 130 131 132 133 134 135 160 161 162 163
+ 164 165 166 167 136 137 138 139 140 141 142 143 168 169 170 171 172 173 174 175
+ Cell_array32x1 $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
