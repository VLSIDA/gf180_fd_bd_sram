* Subcircuit definition of cell ICV_22
.SUBCKT ICV_22 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58
** N=58 EP=58 IP=68 FDC=352
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 27 28
+ 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ ICV_21 $T=-12000 0 0 0 $X=-21340 $Y=-340
X1 1 2 3 4 5 6 7 8 9 10 19 20 21 22 23 24 25 26 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57 58
+ ICV_21 $T=0 0 0 0 $X=-9340 $Y=-340
.ENDS
