* Subcircuit definition of cell din
.SUBCKT din vss 2 3 4 d db 7 8 9 10 11 12 vdd datain men wep
** N=69 EP=16 IP=73 FDC=24
M0 2 4 vss vss nfet_05v0 L=6e-07 W=1.361e-05 AD=5.9884e-12 AS=5.9884e-12 PD=2.81e-05 PS=2.81e-05 NRD=0.0323292 NRS=0.0323292 m=1 nf=1 $X=260 $Y=10430 $D=2
M1 3 wep vss vss nfet_05v0 L=6e-07 W=1.14e-06 AD=7.866e-13 AS=7.923e-13 PD=3.66e-06 PS=3.67e-06 NRD=0.605263 NRS=0.609649 m=1 nf=1 $X=3600 $Y=38320 $D=2
M2 vss 10 4 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=11165 $Y=8655 $D=2
M3 3 wep vdd vdd pfet_05v0 L=6e-07 W=2.97e-06 AD=1.13602e-12 AS=1.7523e-12 PD=4.5e-06 PS=8.3e-06 NRD=0.515152 NRS=0.794613 m=1 nf=2 $X=3025 $Y=35440 $D=8
M4 vdd 2 7 vdd pfet_05v0 L=6e-07 W=1.134e-05 AD=4.9896e-12 AS=4.9896e-12 PD=2.356e-05 PS=2.356e-05 NRD=0.0388007 NRS=0.0388007 m=1 nf=1 $X=6980 $Y=26220 $D=8
X5 4 vdd 10 vdd pfet_05v0_I09 $T=11165 455 0 0 $X=10125 $Y=-165
X6 d 2 3 vdd pmos_1p2$$46889004 $T=2655 26220 0 0 $X=1225 $Y=25510
X7 db 7 3 vdd pmos_1p2$$46889004 $T=4895 26220 0 0 $X=3465 $Y=25510
X9 vdd 2 4 pmos_1p2$$46887980 $T=415 26220 0 0 $X=-1015 $Y=25510
X10 vdd 12 men pmos_1p2$$46273580 $T=2920 7175 1 0 $X=1490 $Y=5355
X11 vdd 11 4 pmos_1p2$$46273580 $T=7060 8140 1 0 $X=5630 $Y=6320
X12 d 2 wep vss nmos_1p2$$46883884 $T=2655 12695 0 0 $X=1510 $Y=12010
X13 db 7 wep vss nmos_1p2$$46883884 $T=4895 12695 0 0 $X=3750 $Y=12010
X14 7 vss 2 vss nmos_1p2$$46883884 $T=7135 12695 0 0 $X=5990 $Y=12010
X15 8 vdd 9 datain 8 vdd pfet_05v0_I03 $T=2765 3195 0 0 $X=1725 $Y=2575
X16 9 10 11 men 12 vdd pfet_05v0_I03 $T=6905 3605 0 0 $X=5865 $Y=2985
X17 8 vss 9 datain 8 vss nfet_05v0_I02 $T=2765 1790 1 0 $X=2085 $Y=210
X18 9 10 11 12 men vss nfet_05v0_I02 $T=6905 725 0 0 $X=6225 $Y=105
X19 vss 12 men vss nmos_1p2$$46563372 $T=3470 9035 0 0 $X=2325 $Y=8350
X20 vss 11 4 vss nmos_1p2$$46563372 $T=7060 10495 1 0 $X=5915 $Y=8860
.ENDS
************* SUBCKT CALLS DEFINITION ***************
.SUBCKT pfet_05v0_I09 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 pfet_05v0 L=6e-07 W=6.81e-06 AD=2.9964e-12 AS=2.9964e-12 PD=1.45e-05 PS=1.45e-05 NRD=0.0646109 NRS=0.0646109 m=1 nf=1 $X=0 $Y=0 $D=8
.ENDS
.SUBCKT pmos_1p2$$46889004 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
X0 1 2 3 4 pfet_05v0_I09 $T=-155 0 0 0 $X=-1195 $Y=-620
.ENDS
.SUBCKT pmos_1p2$$46887980 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=1.361e-05 AD=5.9884e-12 AS=5.9884e-12 PD=2.81e-05 PS=2.81e-05 NRD=0.0323292 NRS=0.0323292 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
.SUBCKT pmos_1p2$$46273580 1 2 3
** N=3 EP=3 IP=3 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=2.28e-06 AD=5.928e-13 AS=1.0032e-12 PD=3.32e-06 PS=6.32e-06 NRD=0.45614 NRS=0.77193 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
.SUBCKT nmos_1p2$$46883884 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nfet_05v0 L=6e-07 W=1.134e-05 AD=4.9896e-12 AS=4.9896e-12 PD=2.356e-05 PS=2.356e-05 NRD=0.0388007 NRS=0.0388007 m=1 nf=1 $X=-155 $Y=0 $D=2
.ENDS
.SUBCKT pfet_05v0_I03 1 2 3 4 5 6
** N=6 EP=6 IP=0 FDC=2
M0 2 4 1 6 pfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=0 $Y=0 $D=8
M1 3 5 2 6 pfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=1120 $Y=0 $D=8
.ENDS
.SUBCKT nfet_05v0_I02 1 2 3 4 5 6
** N=6 EP=6 IP=0 FDC=2
M0 2 4 1 6 nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=0 $Y=0 $D=2
M1 3 5 2 6 nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=1120 $Y=0 $D=2
.ENDS
.SUBCKT nmos_1p2$$46563372 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
M0 2 3 1 4 nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=-155 $Y=0 $D=2
.ENDS
