* Subcircuit definition of cell pmos_1p2$$48624684
.SUBCKT pmos_1p2$$48624684
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
