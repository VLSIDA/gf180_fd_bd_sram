* Subcircuit definition of cell sacntl_2
.SUBCKT sacntl_2 vss 2 pcb 4 5 6 7 8 9 10 11 18 19 20 21 22 23 24 25 26
+ se vdd men
** N=54 EP=23 IP=83 FDC=39
M0 2 11 vss vss nfet_05v0 L=6e-07 W=2.28e-06 AD=5.928e-13 AS=1.0032e-12 PD=3.32e-06 PS=6.32e-06 NRD=0.45614 NRS=0.77193 m=1 nf=2 $X=795 $Y=26115 $D=2
M1 4 men vss vss nfet_05v0 L=6e-07 W=5.7e-06 AD=1.6872e-12 AS=1.6872e-12 PD=9.8e-06 PS=9.8e-06 NRD=1.29825 NRS=1.29825 m=1 nf=5 $X=855 $Y=4275 $D=2
M2 vss 10 pcb vss nfet_05v0 L=6e-07 W=1.589e-05 AD=4.54e-12 AS=4.54e-12 PD=2.216e-05 PS=2.216e-05 NRD=0.881057 NRS=0.881057 m=1 nf=7 $X=1950 $Y=9235 $D=2
M3 5 4 vss vss nfet_05v0 L=6e-07 W=2.86e-06 AD=7.436e-13 AS=1.2584e-12 PD=3.38e-06 PS=6.6e-06 NRD=0.0909091 NRS=0.153846 m=1 nf=1 $X=10910 $Y=8645 $D=2
M4 6 11 5 vss nfet_05v0 L=6e-07 W=2.86e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12030 $Y=8645 $D=2
M5 7 19 6 vss nfet_05v0 L=6e-07 W=2.86e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=13150 $Y=8645 $D=2
M6 8 19 7 vss nfet_05v0 L=6e-07 W=2.86e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=14270 $Y=8645 $D=2
M7 9 11 8 vss nfet_05v0 L=6e-07 W=2.86e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=15390 $Y=8645 $D=2
M8 vss 4 9 vss nfet_05v0 L=6e-07 W=2.86e-06 AD=1.2584e-12 AS=7.436e-13 PD=6.6e-06 PS=3.38e-06 NRD=0.153846 NRS=0.0909091 m=1 nf=1 $X=16510 $Y=8645 $D=2
M9 10 7 vss vss nfet_05v0 L=6e-07 W=5.22e-06 AD=1.3572e-12 AS=2.2968e-12 PD=6.26e-06 PS=1.22e-05 NRD=0.199234 NRS=0.337165 m=1 nf=2 $X=18750 $Y=8895 $D=2
M10 11 20 vss vss nfet_05v0 L=6e-07 W=1.44e-06 AD=6.336e-13 AS=6.336e-13 PD=3.76e-06 PS=3.76e-06 NRD=0.305556 NRS=0.305556 m=1 nf=1 $X=21255 $Y=4090 $D=2
M11 se 19 vss vss nfet_05v0 L=6e-07 W=9.08e-06 AD=2.3608e-12 AS=3.178e-12 PD=1.116e-05 PS=1.642e-05 NRD=0.45815 NRS=0.61674 m=1 nf=4 $X=19460 $Y=25030 $D=2
M12 2 11 vdd vdd pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=3.0008e-12 PD=7.86e-06 PS=1.54e-05 NRD=0.152493 NRS=0.258065 m=1 nf=2 $X=795 $Y=20945 $D=8
M13 4 men vdd vdd pfet_05v0 L=6e-07 W=1.135e-05 AD=3.3596e-12 AS=3.3596e-12 PD=1.658e-05 PS=1.658e-05 NRD=0.651982 NRS=0.651982 m=1 nf=5 $X=855 $Y=590 $D=8
M14 19 2 vdd vdd pfet_05v0 L=6e-07 W=6.81e-06 AD=1.7706e-12 AS=2.1792e-12 PD=8.37e-06 PS=1.1e-05 NRD=0.343612 NRS=0.422907 m=1 nf=3 $X=5370 $Y=20990 $D=8
M15 vdd 4 19 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=8730 $Y=20990 $D=8
M16 pcb 10 vdd vdd pfet_05v0 L=6e-07 W=4.09e-05 AD=1.0634e-11 AS=1.21023e-11 PD=4.61e-05 PS=4.6818e-05 NRD=0.635697 NRS=0.723472 m=1 nf=10 $X=830 $Y=14055 $D=8
M17 7 19 vdd vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.06e-06 PS=9.96e-06 NRD=0.0572687 NRS=0.0969163 m=1 nf=1 $X=14270 $Y=13710 $D=8
M18 vdd 11 7 vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=15390 $Y=13710 $D=8
M19 7 4 vdd vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.9976e-12 AS=1.1804e-12 PD=9.96e-06 PS=5.06e-06 NRD=0.0969163 NRS=0.0572687 m=1 nf=1 $X=16510 $Y=13710 $D=8
M20 vdd 25 26 vdd pfet_05v0 L=6e-07 W=1.2e-06 AD=5.28e-13 AS=5.28e-13 PD=3.28e-06 PS=3.28e-06 NRD=0.366667 NRS=0.366667 m=1 nf=1 $X=18950 $Y=1670 $D=8
M21 10 7 vdd vdd pfet_05v0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=4.3584e-12 PD=2.008e-05 PS=2.008e-05 NRD=0.211454 NRS=0.211454 m=1 nf=3 $X=18750 $Y=13710 $D=8
M22 se 19 vdd vdd pfet_05v0 L=6e-07 W=2.72e-05 AD=7.072e-12 AS=8.0512e-12 PD=3.24e-05 PS=3.856e-05 NRD=0.955882 NRS=1.08824 m=1 nf=10 $X=12740 $Y=20450 $D=8
X23 vdd 11 20 pfet_05v0_I15 $T=21255 985 0 0 $X=20215 $Y=365
X27 vss 18 2 vss nfet_05v0_I10 $T=5370 25030 0 0 $X=4690 $Y=24410
X28 19 18 4 vss nfet_05v0_I10 $T=12415 25030 0 0 $X=11735 $Y=24410
X29 20 vdd 21 4 vss pfet_05v0_I16 $T=8080 1480 0 0 $X=7040 $Y=860
X30 22 vdd 23 21 22 pfet_05v0_I16 $T=11705 1480 0 0 $X=10665 $Y=860
X31 24 vdd 25 23 24 pfet_05v0_I16 $T=15325 1480 0 0 $X=14285 $Y=860
X32 20 vss 21 4 vss nfet_05v0_I17 $T=8080 4420 0 0 $X=7400 $Y=3800
X33 22 vss 23 21 22 nfet_05v0_I17 $T=11705 4420 0 0 $X=11025 $Y=3800
X34 24 vss 25 23 24 nfet_05v0_I17 $T=15325 4420 0 0 $X=14645 $Y=3800
X39 26 vss 25 vss nfet_05v0_I08 $T=18950 4420 0 0 $X=18270 $Y=3800
.ENDS
