* Subcircuit definition of cell ICV_4
.SUBCKT ICV_4 1 2 3 4 14 16 18 19
** N=23 EP=8 IP=30 FDC=40
*.SEEDPROM
M0 1 3 20 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=3180 $Y=16970 $D=2
M1 22 3 1 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=3180 $Y=18260 $D=2
M2 3 4 20 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=3630 $Y=15340 $D=2
M3 3 4 22 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=3630 $Y=19710 $D=2
M4 21 3 3 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=4770 $Y=15340 $D=2
M5 23 3 3 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=4770 $Y=19710 $D=2
M6 2 3 21 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=5220 $Y=16970 $D=2
M7 23 3 2 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=5220 $Y=18260 $D=2
X8 1 2 3 4 14 16 20 21 ICV_3 $T=0 0 0 0 $X=-340 $Y=-340
X9 1 2 3 4 22 23 18 19 ICV_3 $T=0 18000 0 0 $X=-340 $Y=17660
.ENDS
