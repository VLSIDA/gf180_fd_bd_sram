* Subcircuit definition of cell ICV_10
.SUBCKT ICV_10
** N=15 EP=0 IP=20 FDC=0
.ENDS
