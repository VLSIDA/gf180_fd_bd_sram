* Subcircuit definition of cell ICV_24
.SUBCKT ICV_24 1 2 4 7 8 9 10
** N=10 EP=7 IP=14 FDC=8
*.SEEDPROM
M0 1 4 7 4 nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=180 $Y=-1030 $D=2
M1 9 4 1 4 nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=180 $Y=260 $D=2
M2 4 8 7 4 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=-2660 $D=2
M3 4 10 9 4 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=1710 $D=2
M4 8 7 4 4 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=-2660 $D=2
M5 10 9 4 4 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=1710 $D=2
M6 2 4 8 4 nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=2220 $Y=-1030 $D=2
M7 10 4 2 4 nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=2220 $Y=260 $D=2
.ENDS
