* Subcircuit definition of cell ICV_7
.SUBCKT ICV_7 1 3 4 5 6 7 8 9 10 11
** N=15 EP=10 IP=18 FDC=8
*.SEEDPROM
X0 5 4 1 6 7 3 018SRAM_cell1_dummy $T=-3000 0 0 0 $X=-3340 $Y=-340
X1 9 8 1 10 11 3 018SRAM_cell1_dummy $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
