* Subcircuit definition of cell wen_v2
.SUBCKT wen_v2 vss 2 vdd wen clk IGWEN GWE
** N=50 EP=7 IP=93 FDC=30
M0 vss wen 29 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=2545 $Y=1065 $D=2
M1 12 wen vss vss nfet_05v0 L=6e-07 W=6e-06 AD=1.92e-12 AS=1.92e-12 PD=9.92e-06 PS=9.92e-06 NRD=0.48 NRS=0.48 m=1 nf=3 $X=1260 $Y=16070 $D=2
M2 32 clk vss vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=3665 $Y=1065 $D=2
M3 2 32 vss vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=5905 $Y=1475 $D=2
M4 30 32 29 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=8440 $Y=545 $D=2
M5 34 2 30 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=10750 $Y=1860 $D=2
M6 vss 35 34 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=11870 $Y=1860 $D=2
M7 vss 30 35 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=14110 $Y=1860 $D=2
M8 16 35 vss vss nfet_05v0 L=6e-07 W=2.4e-06 AD=6.24e-13 AS=1.056e-12 PD=3.44e-06 PS=6.56e-06 NRD=0.433333 NRS=0.733333 m=1 nf=2 $X=16465 $Y=1620 $D=2
M9 16 2 31 vss nfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=19750 $Y=545 $D=2
M10 33 32 31 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=23090 $Y=1240 $D=2
M11 vss 20 33 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=24210 $Y=1240 $D=2
M12 20 31 vss vss nfet_05v0 L=6e-07 W=6.23e-06 AD=1.78e-12 AS=1.78e-12 PD=1.112e-05 PS=1.112e-05 NRD=2.24719 NRS=2.24719 m=1 nf=7 $X=26535 $Y=1905 $D=2
M13 vdd wen 29 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=2545 $Y=4215 $D=8
M14 32 clk vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=3665 $Y=4215 $D=8
M15 2 32 vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=5905 $Y=4215 $D=8
M16 12 wen vdd vdd pfet_05v0 L=6e-07 W=1.488e-05 AD=3.8688e-12 AS=4.7616e-12 PD=1.8e-05 PS=2.368e-05 NRD=0.629032 NRS=0.774194 m=1 nf=6 $X=1260 $Y=9420 $D=8
M17 30 2 29 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=1.17422e-12 AS=9.988e-13 PD=4.793e-06 PS=5.42e-06 NRD=0.227875 NRS=0.193833 m=1 nf=1 $X=8440 $Y=4215 $D=8
M18 34 32 30 vdd pfet_05v0 L=6e-07 W=9.6e-07 AD=-6.91897e-13 AS=-6.43897e-13 PD=-2.79573e-06 PS=-2.69573e-06 NRD=-0.750757 NRS=-0.698673 m=1 nf=1 $X=10180 $Y=4215 $D=8
M19 vdd 35 34 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=1.14048e-12 PD=5.42e-06 PS=4.72272e-06 NRD=0.193833 NRS=0.221328 m=1 nf=1 $X=11870 $Y=4215 $D=8
M20 vdd 30 35 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=14110 $Y=4215 $D=8
M21 16 35 vdd vdd pfet_05v0 L=6e-07 W=5.68e-06 AD=1.4768e-12 AS=2.4992e-12 PD=6.72e-06 PS=1.312e-05 NRD=0.183099 NRS=0.309859 m=1 nf=2 $X=16465 $Y=4215 $D=8
M22 16 32 31 vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=2.13253e-12 PD=5.58e-06 PS=1.01287e-05 NRD=0.229075 NRS=0.413851 m=1 nf=2 $X=19750 $Y=4215 $D=8
M23 33 2 31 vdd pfet_05v0 L=6e-07 W=9.6e-07 AD=-6.59976e-13 AS=-6.40776e-13 PD=-2.72923e-06 PS=-2.68923e-06 NRD=-0.71612 NRS=-0.695287 m=1 nf=1 $X=22550 $Y=5525 $D=8
M24 vdd 20 33 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=1.12024e-12 PD=5.42e-06 PS=4.68056e-06 NRD=0.193833 NRS=0.2174 m=1 nf=1 $X=24210 $Y=4215 $D=8
M25 20 31 vdd vdd pfet_05v0 L=6e-07 W=1.54e-05 AD=4.4e-12 AS=4.4e-12 PD=2.16e-05 PS=2.16e-05 NRD=0.909091 NRS=0.909091 m=1 nf=7 $X=26535 $Y=4215 $D=8
X48 vss IGWEN 12 nfet_05v0_I08 $T=10115 16070 0 0 $X=9435 $Y=15450
X49 vss GWE 20 nfet_05v0_I08 $T=23345 16070 0 0 $X=22665 $Y=15450
X50 vdd IGWEN 12 pfet_05v0_I06 $T=10115 9420 0 0 $X=9075 $Y=8800
X51 vdd GWE 20 pfet_05v0_I06 $T=23345 9420 0 0 $X=22305 $Y=8800
.ENDS
