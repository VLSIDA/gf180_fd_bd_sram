* Subcircuit definition of cell alatch
.SUBCKT alatch vss ab a vdd enb en
** N=16 EP=6 IP=24 FDC=8
M0 ab 11 vss vss nfet_05v0 L=6e-07 W=3.64e-06 AD=9.464e-13 AS=1.6016e-12 PD=4.68e-06 PS=9.04e-06 NRD=0.285714 NRS=0.483516 m=1 nf=2 $X=2590 $Y=1475 $D=2
M1 vss ab 12 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=3710 $Y=12935 $D=2
M2 a en 11 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=6280 $Y=1020 $D=2
M3 12 enb 11 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=6280 $Y=12935 $D=2
M4 ab 11 vdd vdd pfet_05v0 L=6e-07 W=9.08e-06 AD=2.3608e-12 AS=3.9952e-12 PD=1.012e-05 PS=1.992e-05 NRD=0.114537 NRS=0.193833 m=1 nf=2 $X=2590 $Y=4695 $D=8
M5 a enb 11 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=6280 $Y=5895 $D=8
X10 12 vdd ab vdd pmos_1p2$$47330348_161 $T=3865 11540 1 0 $X=2435 $Y=9910
X11 11 12 en vdd pmos_1p2$$47330348_161 $T=6435 11540 1 0 $X=5005 $Y=9910
.ENDS
