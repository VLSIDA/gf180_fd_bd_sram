* Subcircuit definition of cell M1_PSUB_I03
.SUBCKT M1_PSUB_I03
** N=2001 EP=0 IP=0 FDC=0
.ENDS
