* Subcircuit definition of cell ICV_18
.SUBCKT ICV_18 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46
+ 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66
+ 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86
+ 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106
+ 107 108 109 110 111 112
** N=112 EP=106 IP=152 FDC=704
*.SEEDPROM
X1 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 49 50
+ 51 52 53 54 55 56 57 58 59 60 61 62 63 64
+ ICV_11 $T=0 0 0 0 $X=-340 $Y=-340
X2 7 8 9 10 11 12 13 14 15 16 25 26 27 28 29 30 31 32 65 66
+ 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ ICV_11 $T=12000 0 0 0 $X=11660 $Y=-340
X3 7 8 9 10 11 12 13 14 15 16 33 34 35 36 37 38 39 40 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96
+ ICV_15 $T=30000 0 1 180 $X=26660 $Y=-340
X4 7 8 9 10 11 12 13 14 15 16 41 42 43 44 45 46 47 48 97 98
+ 99 100 101 102 103 104 105 106 107 108 109 110 111 112
+ ICV_15 $T=42000 0 1 180 $X=38660 $Y=-340
.ENDS
