* Subcircuit definition of cell xpredec1_xa
.SUBCKT xpredec1_xa
** N=29 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
