* Subcircuit definition of cell ICV_30
.SUBCKT ICV_30 1 2 3 4 9 11 14 16
** N=16 EP=8 IP=24 FDC=20
*.SEEDPROM
M0 1 12 10 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=8060 $D=8
M1 1 15 13 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=9340 $D=8
M2 12 10 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=8060 $D=8
M3 15 13 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=9340 $D=8
X4 3 4 2 2 2 9 11 10 12 018SRAM_cell1_2x $T=0 0 0 0 $X=-340 $Y=-340
X5 3 4 2 2 2 13 15 14 16 018SRAM_cell1_2x $T=0 9000 0 0 $X=-340 $Y=8660
.ENDS
