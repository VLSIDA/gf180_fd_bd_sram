* Subcircuit definition of cell ICV_5
.SUBCKT ICV_5 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19
** N=27 EP=18 IP=30 FDC=16
*.SEEDPROM
X0 1 3 4 5 6 7 8 9 10 11 ICV_4 $T=-6000 0 0 0 $X=-9340 $Y=-340
X1 1 3 12 13 14 15 16 17 18 19 ICV_4 $T=0 0 0 0 $X=-3340 $Y=-340
.ENDS
