* Subcircuit definition of cell ICV_14
.SUBCKT ICV_14 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
** N=29 EP=17 IP=32 FDC=16
*.SEEDPROM
X0 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 ICV_13 $T=-3000 0 0 0 $X=-12340 $Y=-340
.ENDS
