* Subcircuit definition of cell ICV_20
.SUBCKT ICV_20 1 2 4 5 7 8
** N=8 EP=6 IP=10 FDC=4
*.SEEDPROM
M0 1 7 4 1 nfet_05v0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=3510 $Y=1700 $D=2
M1 8 5 1 1 nfet_05v0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=6870 $Y=1700 $D=2
M2 2 7 4 2 pfet_05v0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=3510 $Y=14855 $D=8
M3 8 5 2 2 pfet_05v0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=6870 $Y=14855 $D=8
.ENDS
