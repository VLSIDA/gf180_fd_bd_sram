* Subcircuit definition of cell nfet_05v0_I10
.SUBCKT nfet_05v0_I10
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
