* Subcircuit definition of cell new_dummyrow_unit
.SUBCKT new_dummyrow_unit 7 9 43 45 47 49 51 53 55 57 59 61 63 65 67 69 71 73 75 77
+ 79 81 83 85 87 89 91 93 95 97 99 101 103 105
** N=105 EP=34 IP=120 FDC=64
*.SEEDPROM
X0 7 9 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 ICV_8 $T=3310 885 1 180 $X=-30 $Y=545
X1 7 9 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 ICV_8 $T=15310 885 1 180 $X=11970 $Y=545
X2 7 9 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 ICV_8 $T=30310 885 1 180 $X=26970 $Y=545
X3 7 9 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 ICV_8 $T=42310 885 1 180 $X=38970 $Y=545
.ENDS
