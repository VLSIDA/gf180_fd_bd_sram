* Subcircuit definition of cell M1_PSUB_I06
.SUBCKT M1_PSUB_I06
** N=1191 EP=0 IP=0 FDC=0
.ENDS
