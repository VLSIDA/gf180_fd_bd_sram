* Subcircuit definition of cell nfet_05v0_I12
.SUBCKT nfet_05v0_I12 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 2 4 1 2 nfet_05v0 L=6e-07 W=6e-07 AD=1.56e-13 AS=2.64e-13 PD=1.12e-06 PS=2.08e-06 NRD=0.433333 NRS=0.733333 m=1 nf=1 $X=0 $Y=0 $D=2
M1 3 5 2 2 nfet_05v0 L=6e-07 W=6e-07 AD=2.64e-13 AS=1.56e-13 PD=2.08e-06 PS=1.12e-06 NRD=0.733333 NRS=0.433333 m=1 nf=1 $X=1120 $Y=0 $D=2
.ENDS
