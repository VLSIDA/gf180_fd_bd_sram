* Subcircuit definition of cell M1_PACTIVE$10
.SUBCKT M1_PACTIVE$10
** N=13 EP=0 IP=0 FDC=0
.ENDS
