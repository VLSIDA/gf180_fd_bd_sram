* Subcircuit definition of cell gf180mcu_fd_ip_sram__sram512x8m8wm1
.SUBCKT gf180mcu_fd_ip_sram__sram512x8m8wm1 A[8] A[7] A[6] A[5] A[4] A[3] A[2]
+ A[1] A[0] CEN CLK D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] GWEN Q[7] Q[6]
+ Q[5] Q[4] Q[3] Q[2] Q[1] Q[0] VDD VSS WEN[7] WEN[6] WEN[5] WEN[4] WEN[3]
+ WEN[2] WEN[1] WEN[0]
** N=24897 EP=38 IP=4916 FDC=29933
M0 23498 VSS 703 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=120390 $Y=176390 $D=2
M1 703 VSS 23500 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=120390 $Y=472100 $D=2
M2 VSS 23497 23498 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=120840 $Y=177840 $D=2
M3 VSS 23499 23500 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=120840 $Y=470470 $D=2
M4 23497 23498 VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=121980 $Y=177840 $D=2
M5 23499 23500 VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=121980 $Y=470470 $D=2
M6 23497 VSS 702 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=122430 $Y=176390 $D=2
M7 702 VSS 23499 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=122430 $Y=472100 $D=2
M8 VSS 24106 23202 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=168355 $Y=180895 $D=2
M9 24106 24042 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=183295 $D=2
M10 VSS 24044 24108 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=213375 $D=2
M11 VSS 24108 23209 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=214655 $D=2
M12 VSS 24110 23210 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=216895 $D=2
M13 24110 24046 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=219295 $D=2
M14 VSS 24048 24112 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=249375 $D=2
M15 VSS 24112 23217 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=250655 $D=2
M16 VSS 24114 23218 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=252895 $D=2
M17 24114 24050 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=255295 $D=2
M18 VSS 24052 24116 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=285375 $D=2
M19 VSS 24116 23225 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=286655 $D=2
M20 VSS 24118 23226 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=288895 $D=2
M21 24118 24054 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=291295 $D=2
M22 VSS 24056 24120 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=321375 $D=2
M23 VSS 24120 23233 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=322655 $D=2
M24 VSS 24122 23234 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=324895 $D=2
M25 24122 24058 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=327295 $D=2
M26 VSS 24060 24124 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=357375 $D=2
M27 VSS 24124 23241 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=358655 $D=2
M28 VSS 24126 23242 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=360895 $D=2
M29 24126 24062 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=363295 $D=2
M30 VSS 24064 24128 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=393375 $D=2
M31 VSS 24128 23249 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=394655 $D=2
M32 VSS 24130 23250 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=396895 $D=2
M33 24130 24066 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=399295 $D=2
M34 VSS 24068 24132 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=429375 $D=2
M35 VSS 24132 23257 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=430655 $D=2
M36 VSS 24134 23258 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=432895 $D=2
M37 24134 24070 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=435295 $D=2
M38 VSS 24072 24136 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=465375 $D=2
M39 VSS 24136 23265 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=168355 $Y=466655 $D=2
M40 24042 24043 VSS VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=198635 $Y=180895 $D=2
M41 VSS 24045 24044 VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=215775 $D=2
M42 24046 24047 VSS VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=216895 $D=2
M43 VSS 24049 24048 VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=251775 $D=2
M44 24050 24051 VSS VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=252895 $D=2
M45 VSS 24053 24052 VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=287775 $D=2
M46 24054 24055 VSS VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=288895 $D=2
M47 VSS 24057 24056 VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=323775 $D=2
M48 24058 24059 VSS VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=324895 $D=2
M49 VSS 24061 24060 VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=359775 $D=2
M50 24062 24063 VSS VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=360895 $D=2
M51 VSS 24065 24064 VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=395775 $D=2
M52 24066 24067 VSS VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=396895 $D=2
M53 VSS 24069 24068 VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=431775 $D=2
M54 24070 24071 VSS VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=432895 $D=2
M55 VSS 24073 24072 VSS nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=198635 $Y=467775 $D=2
M56 2 VDD 1 VSS nfet_05v0 L=6e-07 W=6.59e-06 AD=2.8996e-12 AS=2.8996e-12 PD=1.406e-05 PS=1.406e-05 NRD=0.0667678 NRS=0.0667678 m=1 nf=1 $X=204815 $Y=471000 $D=2
M57 24707 1040 VSS VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=7.32375e-13 AS=2.079e-12 PD=3.615e-06 PS=7.62e-06 NRD=0.0738095 NRS=0.209524 m=1 nf=1 $X=218475 $Y=180950 $D=2
M58 24706 1044 24707 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=182015 $D=2
M59 24043 1052 24706 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=183135 $D=2
M60 24708 1045 24045 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=213535 $D=2
M61 24709 1044 24708 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=214655 $D=2
M62 VSS 1040 24709 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=215720 $D=2
M63 24711 1040 VSS VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=216950 $D=2
M64 24710 1043 24711 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=218015 $D=2
M65 24047 1052 24710 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=219135 $D=2
M66 24712 1045 24049 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=249535 $D=2
M67 24713 1043 24712 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=250655 $D=2
M68 VSS 1040 24713 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=251720 $D=2
M69 24715 1040 VSS VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=252950 $D=2
M70 24714 1042 24715 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=254015 $D=2
M71 24051 1052 24714 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=255135 $D=2
M72 24716 1045 24053 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=285535 $D=2
M73 24717 1042 24716 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=286655 $D=2
M74 VSS 1040 24717 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=287720 $D=2
M75 24719 1040 VSS VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=288950 $D=2
M76 24718 1041 24719 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=290015 $D=2
M77 24055 1052 24718 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=291135 $D=2
M78 24720 1045 24057 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=321535 $D=2
M79 24721 1041 24720 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=322655 $D=2
M80 VSS 1040 24721 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=323720 $D=2
M81 24723 1038 VSS VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=324950 $D=2
M82 24722 1044 24723 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=326015 $D=2
M83 24059 1052 24722 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=327135 $D=2
M84 24724 1045 24061 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=357535 $D=2
M85 24725 1044 24724 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=358655 $D=2
M86 VSS 1038 24725 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=359720 $D=2
M87 24727 1038 VSS VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=360950 $D=2
M88 24726 1043 24727 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=362015 $D=2
M89 24063 1052 24726 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=363135 $D=2
M90 24728 1045 24065 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=393535 $D=2
M91 24729 1043 24728 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=394655 $D=2
M92 VSS 1038 24729 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=395720 $D=2
M93 24731 1038 VSS VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=396950 $D=2
M94 24730 1042 24731 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=398015 $D=2
M95 24067 1052 24730 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=399135 $D=2
M96 24732 1045 24069 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=429535 $D=2
M97 24733 1042 24732 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=430655 $D=2
M98 VSS 1038 24733 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=431720 $D=2
M99 24735 1038 VSS VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=432950 $D=2
M100 24734 1041 24735 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=434015 $D=2
M101 24071 1052 24734 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=435135 $D=2
M102 24736 1045 24073 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=465535 $D=2
M103 24737 1041 24736 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=466655 $D=2
M104 VSS 1038 24737 VSS nfet_05v0 L=6e-07 W=3.15e-06 AD=2.079e-12 AS=7.32375e-13 PD=7.62e-06 PS=3.615e-06 NRD=0.209524 NRS=0.0738095 m=1 nf=1 $X=218475 $Y=467720 $D=2
M105 VSS 1 1000 VSS nfet_05v0 L=6e-07 W=1.36e-06 AD=3.536e-13 AS=5.984e-13 PD=1.88e-06 PS=3.6e-06 NRD=0.191176 NRS=0.323529 m=1 nf=1 $X=233770 $Y=54135 $D=2
M106 1000 CLK VSS VSS nfet_05v0 L=6e-07 W=1.36e-06 AD=5.984e-13 AS=3.536e-13 PD=3.6e-06 PS=1.88e-06 NRD=0.323529 NRS=0.191176 m=1 nf=1 $X=234890 $Y=54135 $D=2
M107 616 619 VSS VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=242235 $Y=54135 $D=2
M108 281 1006 VSS VSS nfet_05v0 L=1e-06 W=6e-07 AD=2.64e-13 AS=2.64e-13 PD=2.08e-06 PS=2.08e-06 NRD=0.733333 NRS=0.733333 m=1 nf=1 $X=243265 $Y=46010 $D=2
M109 CEN 1000 619 VSS nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=245925 $Y=54135 $D=2
M110 250 468 VSS VSS nfet_05v0 L=6e-07 W=4.99e-05 AD=1.47704e-11 AS=1.47704e-11 PD=6.284e-05 PS=6.284e-05 NRD=0.148297 NRS=0.148297 m=1 nf=5 $X=241995 $Y=72320 $D=2
M111 317 281 VSS VSS nfet_05v0 L=6e-07 W=7.5e-07 AD=3.3e-13 AS=3.3e-13 PD=2.38e-06 PS=2.38e-06 NRD=0.586667 NRS=0.586667 m=1 nf=1 $X=246495 $Y=46075 $D=2
M112 354 317 VSS VSS nfet_05v0 L=6e-07 W=3.02e-06 AD=1.3288e-12 AS=1.3288e-12 PD=6.92e-06 PS=6.92e-06 NRD=0.145695 NRS=0.145695 m=1 nf=1 $X=249065 $Y=46070 $D=2
M113 24027 354 VSS VSS nfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=1.34946e-11 PD=2.32e-05 PS=4.655e-05 NRD=0.0114638 NRS=0.0262346 m=1 nf=1 $X=256125 $Y=28435 $D=2
M114 VSS 24107 23266 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=252270 $Y=180895 $D=2
M115 24107 24042 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=183295 $D=2
M116 VSS 24044 24109 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=213375 $D=2
M117 VSS 24109 23273 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=214655 $D=2
M118 VSS 24111 23274 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=216895 $D=2
M119 24111 24046 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=219295 $D=2
M120 VSS 24048 24113 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=249375 $D=2
M121 VSS 24113 23281 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=250655 $D=2
M122 VSS 24115 23282 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=252895 $D=2
M123 24115 24050 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=255295 $D=2
M124 VSS 24052 24117 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=285375 $D=2
M125 VSS 24117 23289 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=286655 $D=2
M126 VSS 24119 23290 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=288895 $D=2
M127 24119 24054 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=291295 $D=2
M128 VSS 24056 24121 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=321375 $D=2
M129 VSS 24121 23297 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=322655 $D=2
M130 VSS 24123 23298 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=324895 $D=2
M131 24123 24058 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=327295 $D=2
M132 VSS 24060 24125 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=357375 $D=2
M133 VSS 24125 23305 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=358655 $D=2
M134 VSS 24127 23306 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=360895 $D=2
M135 24127 24062 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=363295 $D=2
M136 VSS 24064 24129 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=393375 $D=2
M137 VSS 24129 23313 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=394655 $D=2
M138 VSS 24131 23314 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=396895 $D=2
M139 24131 24066 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=399295 $D=2
M140 VSS 24068 24133 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=429375 $D=2
M141 VSS 24133 23321 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=430655 $D=2
M142 VSS 24135 23322 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=432895 $D=2
M143 24135 24070 VSS VSS nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=435295 $D=2
M144 VSS 24072 24137 VSS nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=465375 $D=2
M145 VSS 24137 23329 VSS nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=252270 $Y=466655 $D=2
M146 24028 CLK 24027 VSS nfet_05v0 L=6e-07 W=2.268e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=257245 $Y=28435 $D=2
M147 445 616 24028 VSS nfet_05v0 L=6e-07 W=2.268e-05 AD=1.33812e-11 AS=5.8968e-12 PD=4.654e-05 PS=2.32e-05 NRD=0.0260141 NRS=0.0114638 m=1 nf=1 $X=258365 $Y=28435 $D=2
M148 24029 495 VSS VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=4.7177e-12 AS=1.07963e-11 PD=1.8665e-05 PS=3.748e-05 NRD=0.014329 NRS=0.0327914 m=1 nf=1 $X=262120 $Y=29545 $D=2
M149 468 445 24029 VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=263240 $Y=29545 $D=2
M150 24030 445 468 VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=264360 $Y=29545 $D=2
M151 VSS 495 24030 VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=1.07055e-11 AS=4.7177e-12 PD=3.747e-05 PS=1.8665e-05 NRD=0.0325158 NRS=0.014329 m=1 nf=1 $X=265480 $Y=29545 $D=2
M152 24031 468 VSS VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=1.16905e-12 AS=2.7013e-12 PD=5.055e-06 PS=1.027e-05 NRD=0.0567181 NRS=0.131057 m=1 nf=1 $X=268545 $Y=43150 $D=2
M153 495 607 24031 VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=2.27e-14 AS=-2.27e-14 PD=1e-08 PS=-1e-08 NRD=0.00110132 NRS=-0.00110132 m=1 nf=1 $X=269660 $Y=43150 $D=2
M154 24032 607 495 VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=-2.27e-14 AS=2.27e-14 PD=-1e-08 PS=1e-08 NRD=-0.00110132 NRS=0.00110132 m=1 nf=1 $X=270785 $Y=43150 $D=2
M155 VSS 468 24032 VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=2.7013e-12 AS=1.16905e-12 PD=1.027e-05 PS=5.055e-06 NRD=0.131057 NRS=0.0567181 m=1 nf=1 $X=271900 $Y=43150 $D=2
M156 1 250 VSS VSS nfet_05v0 L=6e-07 W=0.0001474 AD=3.8324e-11 AS=4.09772e-11 PD=0.0001578 PS=0.00017326 NRD=0.705563 NRS=0.75441 m=1 nf=20 $X=253180 $Y=76320 $D=2
M157 23502 VSS 705 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=304270 $Y=176390 $D=2
M158 705 VSS 23504 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=304270 $Y=472100 $D=2
M159 VSS 23501 23502 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=304720 $Y=177840 $D=2
M160 VSS 23503 23504 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=304720 $Y=470470 $D=2
M161 23501 23502 VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=305860 $Y=177840 $D=2
M162 23503 23504 VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=305860 $Y=470470 $D=2
M163 23501 VSS 704 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=306310 $Y=176390 $D=2
M164 704 VSS 23503 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=306310 $Y=472100 $D=2
M165 24074 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=418270 $Y=176390 $D=2
M166 614 VSS 24076 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=211100 $D=2
M167 24078 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=212390 $D=2
M168 614 VSS 24080 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=247100 $D=2
M169 24082 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=248390 $D=2
M170 614 VSS 24084 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=283100 $D=2
M171 24086 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=284390 $D=2
M172 614 VSS 24088 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=319100 $D=2
M173 24090 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=320390 $D=2
M174 614 VSS 24092 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=355100 $D=2
M175 24094 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=356390 $D=2
M176 614 VSS 24096 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=391100 $D=2
M177 24098 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=392390 $D=2
M178 614 VSS 24100 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=427100 $D=2
M179 24102 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=428390 $D=2
M180 614 1002 24104 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=463100 $D=2
M181 23859 1002 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=464390 $D=2
M182 614 1002 23857 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=418270 $Y=472100 $D=2
M183 VSS VDD 24074 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=177840 $D=2
M184 VSS VDD 24076 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=209470 $D=2
M185 VSS VDD 24078 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=213840 $D=2
M186 VSS VDD 24080 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=245470 $D=2
M187 VSS VDD 24082 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=249840 $D=2
M188 VSS VDD 24084 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=281470 $D=2
M189 VSS VDD 24086 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=285840 $D=2
M190 VSS VDD 24088 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=317470 $D=2
M191 VSS VDD 24090 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=321840 $D=2
M192 VSS VDD 24092 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=353470 $D=2
M193 VSS VDD 24094 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=357840 $D=2
M194 VSS VDD 24096 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=389470 $D=2
M195 VSS VDD 24098 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=393840 $D=2
M196 VSS VDD 24100 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=425470 $D=2
M197 VSS VDD 24102 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=429840 $D=2
M198 VSS VDD 24104 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=461470 $D=2
M199 VSS VDD 23859 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=465840 $D=2
M200 VSS VDD 23857 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=470470 $D=2
M201 24075 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=177840 $D=2
M202 24077 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=209470 $D=2
M203 24079 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=213840 $D=2
M204 24081 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=245470 $D=2
M205 24083 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=249840 $D=2
M206 24085 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=281470 $D=2
M207 24087 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=285840 $D=2
M208 24089 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=317470 $D=2
M209 24091 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=321840 $D=2
M210 24093 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=353470 $D=2
M211 24095 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=357840 $D=2
M212 24097 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=389470 $D=2
M213 24099 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=393840 $D=2
M214 24101 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=425470 $D=2
M215 24103 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=429840 $D=2
M216 24105 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=461470 $D=2
M217 23860 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=465840 $D=2
M218 23858 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=470470 $D=2
M219 606 614 VSS VSS nfet_05v0 L=6e-07 W=2.76e-06 AD=7.176e-13 AS=1.2144e-12 PD=3.8e-06 PS=7.28e-06 NRD=0.376812 NRS=0.637681 m=1 nf=2 $X=418770 $Y=94540 $D=2
M220 607 606 VSS VSS nfet_05v0 L=6e-07 W=1.7e-05 AD=4.42e-12 AS=7.48e-12 PD=1.804e-05 PS=3.576e-05 NRD=0.0611765 NRS=0.103529 m=1 nf=2 $X=418790 $Y=79115 $D=2
M221 613 VDD VSS VSS nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=5.016e-13 PD=2.18e-06 PS=4.04e-06 NRD=0.912281 NRS=1.54386 m=1 nf=2 $X=419015 $Y=110805 $D=2
M222 24075 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=420310 $Y=176390 $D=2
M223 615 VSS 24077 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=211100 $D=2
M224 24079 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=212390 $D=2
M225 615 VSS 24081 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=247100 $D=2
M226 24083 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=248390 $D=2
M227 615 VSS 24085 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=283100 $D=2
M228 24087 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=284390 $D=2
M229 615 VSS 24089 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=319100 $D=2
M230 24091 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=320390 $D=2
M231 615 VSS 24093 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=355100 $D=2
M232 24095 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=356390 $D=2
M233 615 VSS 24097 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=391100 $D=2
M234 24099 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=392390 $D=2
M235 615 VSS 24101 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=427100 $D=2
M236 24103 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=428390 $D=2
M237 615 1002 24105 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=463100 $D=2
M238 23860 1002 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=464390 $D=2
M239 615 1002 23858 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=420310 $Y=472100 $D=2
M240 VDD 23446 23448 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=179690 $D=8
M241 VDD 24167 24166 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=180970 $D=8
M242 VDD 24175 24174 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=323690 $D=8
M243 VDD 24183 24182 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=324970 $D=8
M244 VDD 24191 24190 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=467690 $D=8
M245 VDD 23534 23536 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=468970 $D=8
M246 23446 23448 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=179690 $D=8
M247 24167 24166 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=180970 $D=8
M248 24175 24174 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=323690 $D=8
M249 24183 24182 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=324970 $D=8
M250 24191 24190 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=467690 $D=8
M251 23534 23536 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=468970 $D=8
M252 23915 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=13620 $Y=160970 $D=8
M253 23916 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=13620 $Y=164845 $D=8
M254 24138 23885 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=13835 $Y=112830 $D=8
M255 VDD 23442 23444 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=179690 $D=8
M256 VDD 24169 24168 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=180970 $D=8
M257 VDD 24177 24176 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=323690 $D=8
M258 VDD 24185 24184 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=324970 $D=8
M259 VDD 24193 24192 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=467690 $D=8
M260 VDD 23530 23532 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=468970 $D=8
M261 23442 23444 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=179690 $D=8
M262 24169 24168 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=180970 $D=8
M263 24177 24176 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=323690 $D=8
M264 24185 24184 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=324970 $D=8
M265 24193 24192 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=467690 $D=8
M266 23530 23532 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=468970 $D=8
M267 24139 23884 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=16365 $Y=112830 $D=8
M268 23918 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=16720 $Y=160970 $D=8
M269 23917 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=16720 $Y=164845 $D=8
M270 VDD 23438 23440 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=179690 $D=8
M271 VDD 24171 24170 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=180970 $D=8
M272 VDD 24179 24178 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=323690 $D=8
M273 VDD 24187 24186 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=324970 $D=8
M274 VDD 24195 24194 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=467690 $D=8
M275 VDD 23526 23528 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=468970 $D=8
M276 23438 23440 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=179690 $D=8
M277 24171 24170 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=180970 $D=8
M278 24179 24178 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=323690 $D=8
M279 24187 24186 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=324970 $D=8
M280 24195 24194 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=467690 $D=8
M281 23526 23528 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=468970 $D=8
M282 23919 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=19815 $Y=160970 $D=8
M283 23920 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=19815 $Y=164845 $D=8
M284 24140 23883 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=20030 $Y=112830 $D=8
M285 VDD 23434 23436 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=179690 $D=8
M286 VDD 24173 24172 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=180970 $D=8
M287 VDD 24181 24180 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=323690 $D=8
M288 VDD 24189 24188 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=324970 $D=8
M289 VDD 24197 24196 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=467690 $D=8
M290 VDD 23522 23524 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=468970 $D=8
M291 23434 23436 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=179690 $D=8
M292 24173 24172 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=180970 $D=8
M293 24181 24180 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=323690 $D=8
M294 24189 24188 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=324970 $D=8
M295 24197 24196 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=467690 $D=8
M296 23522 23524 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=468970 $D=8
M297 24141 23882 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=22560 $Y=112830 $D=8
M298 23922 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=22915 $Y=160970 $D=8
M299 23921 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=22915 $Y=164845 $D=8
M300 VDD 23342 23344 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=179690 $D=8
M301 VDD 24263 24262 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=180970 $D=8
M302 VDD 24287 24286 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=323690 $D=8
M303 VDD 24311 24310 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=324970 $D=8
M304 VDD 24335 24334 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=467690 $D=8
M305 VDD 23518 23520 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=468970 $D=8
M306 23342 23344 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=179690 $D=8
M307 24263 24262 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=180970 $D=8
M308 24287 24286 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=323690 $D=8
M309 24311 24310 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=324970 $D=8
M310 24335 24334 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=467690 $D=8
M311 23518 23520 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=468970 $D=8
M312 23923 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=26005 $Y=160970 $D=8
M313 23924 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=26005 $Y=164845 $D=8
M314 24142 23881 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=26220 $Y=112830 $D=8
M315 VDD 23338 23340 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=179690 $D=8
M316 VDD 24265 24264 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=180970 $D=8
M317 VDD 24289 24288 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=323690 $D=8
M318 VDD 24313 24312 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=324970 $D=8
M319 VDD 24337 24336 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=467690 $D=8
M320 VDD 23514 23516 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=468970 $D=8
M321 23338 23340 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=179690 $D=8
M322 24265 24264 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=180970 $D=8
M323 24289 24288 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=323690 $D=8
M324 24313 24312 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=324970 $D=8
M325 24337 24336 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=467690 $D=8
M326 23514 23516 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=468970 $D=8
M327 24143 23880 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=28750 $Y=112830 $D=8
M328 23926 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=29105 $Y=160970 $D=8
M329 23925 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=29105 $Y=164845 $D=8
M330 VDD 23350 23352 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=179690 $D=8
M331 VDD 24267 24266 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=180970 $D=8
M332 VDD 24291 24290 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=323690 $D=8
M333 VDD 24315 24314 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=324970 $D=8
M334 VDD 24339 24338 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=467690 $D=8
M335 VDD 23510 23512 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=468970 $D=8
M336 23350 23352 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=179690 $D=8
M337 24267 24266 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=180970 $D=8
M338 24291 24290 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=323690 $D=8
M339 24315 24314 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=324970 $D=8
M340 24339 24338 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=467690 $D=8
M341 23510 23512 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=468970 $D=8
M342 23927 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=32200 $Y=160970 $D=8
M343 23928 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=32200 $Y=164845 $D=8
M344 24144 23879 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=32415 $Y=112830 $D=8
M345 VDD 23346 23348 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=179690 $D=8
M346 VDD 24269 24268 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=180970 $D=8
M347 VDD 24293 24292 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=323690 $D=8
M348 VDD 24317 24316 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=324970 $D=8
M349 VDD 24341 24340 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=467690 $D=8
M350 VDD 23506 23508 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=468970 $D=8
M351 23346 23348 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=179690 $D=8
M352 24269 24268 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=180970 $D=8
M353 24293 24292 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=323690 $D=8
M354 24317 24316 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=324970 $D=8
M355 24341 24340 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=467690 $D=8
M356 23506 23508 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=468970 $D=8
M357 24034 23878 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=34945 $Y=112830 $D=8
M358 1064 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=35120 $Y=160970 $D=8
M359 1065 23198 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=35120 $Y=164845 $D=8
M360 1076 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=38575 $Y=160970 $D=8
M361 1077 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=38575 $Y=164845 $D=8
M362 VDD 23566 23568 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=179690 $D=8
M363 VDD 24284 24285 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=180970 $D=8
M364 VDD 24308 24309 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=323690 $D=8
M365 VDD 24332 24333 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=324970 $D=8
M366 VDD 24356 24357 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=467690 $D=8
M367 VDD 23598 23600 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=468970 $D=8
M368 24038 23885 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=38620 $Y=112830 $D=8
M369 23566 23568 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=179690 $D=8
M370 24284 24285 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=180970 $D=8
M371 24308 24309 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=323690 $D=8
M372 24332 24333 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=324970 $D=8
M373 24356 24357 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=467690 $D=8
M374 23598 23600 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=468970 $D=8
M375 24652 23884 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=41145 $Y=112830 $D=8
M376 23983 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=41500 $Y=160970 $D=8
M377 23984 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=41500 $Y=164845 $D=8
M378 VDD 23562 23564 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=179690 $D=8
M379 VDD 24282 24283 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=180970 $D=8
M380 VDD 24306 24307 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=323690 $D=8
M381 VDD 24330 24331 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=324970 $D=8
M382 VDD 24354 24355 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=467690 $D=8
M383 VDD 23594 23596 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=468970 $D=8
M384 23562 23564 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=179690 $D=8
M385 24282 24283 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=180970 $D=8
M386 24306 24307 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=323690 $D=8
M387 24330 24331 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=324970 $D=8
M388 24354 24355 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=467690 $D=8
M389 23594 23596 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=468970 $D=8
M390 23982 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=44595 $Y=160970 $D=8
M391 23981 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=44595 $Y=164845 $D=8
M392 VDD 23558 23560 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=179690 $D=8
M393 VDD 24280 24281 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=180970 $D=8
M394 VDD 24304 24305 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=323690 $D=8
M395 VDD 24328 24329 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=324970 $D=8
M396 VDD 24352 24353 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=467690 $D=8
M397 VDD 23590 23592 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=468970 $D=8
M398 24651 23883 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=44810 $Y=112830 $D=8
M399 23558 23560 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=179690 $D=8
M400 24280 24281 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=180970 $D=8
M401 24304 24305 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=323690 $D=8
M402 24328 24329 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=324970 $D=8
M403 24352 24353 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=467690 $D=8
M404 23590 23592 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=468970 $D=8
M405 24650 23882 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=47340 $Y=112830 $D=8
M406 23979 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=47695 $Y=160970 $D=8
M407 23980 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=47695 $Y=164845 $D=8
M408 VDD 23554 23556 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=179690 $D=8
M409 VDD 24278 24279 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=180970 $D=8
M410 VDD 24302 24303 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=323690 $D=8
M411 VDD 24326 24327 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=324970 $D=8
M412 VDD 24350 24351 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=467690 $D=8
M413 VDD 23586 23588 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=468970 $D=8
M414 23554 23556 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=179690 $D=8
M415 24278 24279 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=180970 $D=8
M416 24302 24303 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=323690 $D=8
M417 24326 24327 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=324970 $D=8
M418 24350 24351 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=467690 $D=8
M419 23586 23588 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=468970 $D=8
M420 VDD 23550 23552 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=179690 $D=8
M421 VDD 24276 24277 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=180970 $D=8
M422 VDD 24300 24301 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=323690 $D=8
M423 VDD 24324 24325 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=324970 $D=8
M424 VDD 24348 24349 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=467690 $D=8
M425 VDD 23582 23584 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=468970 $D=8
M426 23978 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=50785 $Y=160970 $D=8
M427 23977 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=50785 $Y=164845 $D=8
M428 24649 23881 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=51000 $Y=112830 $D=8
M429 23550 23552 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=179690 $D=8
M430 24276 24277 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=180970 $D=8
M431 24300 24301 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=323690 $D=8
M432 24324 24325 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=324970 $D=8
M433 24348 24349 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=467690 $D=8
M434 23582 23584 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=468970 $D=8
M435 24648 23880 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=53530 $Y=112830 $D=8
M436 VDD 23546 23548 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=179690 $D=8
M437 VDD 24274 24275 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=180970 $D=8
M438 VDD 24298 24299 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=323690 $D=8
M439 VDD 24322 24323 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=324970 $D=8
M440 VDD 24346 24347 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=467690 $D=8
M441 VDD 23578 23580 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=468970 $D=8
M442 23975 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=53885 $Y=160970 $D=8
M443 23976 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=53885 $Y=164845 $D=8
M444 23546 23548 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=179690 $D=8
M445 24274 24275 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=180970 $D=8
M446 24298 24299 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=323690 $D=8
M447 24322 24323 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=324970 $D=8
M448 24346 24347 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=467690 $D=8
M449 23578 23580 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=468970 $D=8
M450 VDD 23542 23544 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=179690 $D=8
M451 VDD 24272 24273 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=180970 $D=8
M452 VDD 24296 24297 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=323690 $D=8
M453 VDD 24320 24321 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=324970 $D=8
M454 VDD 24344 24345 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=467690 $D=8
M455 VDD 23574 23576 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=468970 $D=8
M456 23974 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=56980 $Y=160970 $D=8
M457 23973 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=56980 $Y=164845 $D=8
M458 24647 23879 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=57195 $Y=112830 $D=8
M459 23542 23544 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=179690 $D=8
M460 24272 24273 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=180970 $D=8
M461 24296 24297 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=323690 $D=8
M462 24320 24321 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=324970 $D=8
M463 24344 24345 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=467690 $D=8
M464 23574 23576 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=468970 $D=8
M465 VDD 23538 23540 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=179690 $D=8
M466 VDD 24270 24271 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=180970 $D=8
M467 VDD 24294 24295 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=323690 $D=8
M468 VDD 24318 24319 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=324970 $D=8
M469 VDD 24342 24343 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=467690 $D=8
M470 VDD 23570 23572 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=468970 $D=8
M471 24646 23878 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=59725 $Y=112830 $D=8
M472 23971 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=60080 $Y=160970 $D=8
M473 23972 1074 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=60080 $Y=164845 $D=8
M474 23538 23540 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=179690 $D=8
M475 24270 24271 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=180970 $D=8
M476 24294 24295 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=323690 $D=8
M477 24318 24319 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=324970 $D=8
M478 24342 24343 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=467690 $D=8
M479 23570 23572 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=468970 $D=8
M480 VDD 23462 23464 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=179690 $D=8
M481 VDD 24199 24198 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=180970 $D=8
M482 VDD 24207 24206 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=323690 $D=8
M483 VDD 24215 24214 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=324970 $D=8
M484 VDD 24223 24222 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=467690 $D=8
M485 VDD 23630 23632 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=468970 $D=8
M486 23462 23464 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=179690 $D=8
M487 24199 24198 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=180970 $D=8
M488 24207 24206 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=323690 $D=8
M489 24215 24214 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=324970 $D=8
M490 24223 24222 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=467690 $D=8
M491 23630 23632 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=468970 $D=8
M492 23929 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=67620 $Y=160970 $D=8
M493 23930 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=67620 $Y=164845 $D=8
M494 24145 23885 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=67835 $Y=112830 $D=8
M495 VDD 23458 23460 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=179690 $D=8
M496 VDD 24201 24200 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=180970 $D=8
M497 VDD 24209 24208 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=323690 $D=8
M498 VDD 24217 24216 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=324970 $D=8
M499 VDD 24225 24224 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=467690 $D=8
M500 VDD 23626 23628 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=468970 $D=8
M501 23458 23460 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=179690 $D=8
M502 24201 24200 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=180970 $D=8
M503 24209 24208 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=323690 $D=8
M504 24217 24216 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=324970 $D=8
M505 24225 24224 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=467690 $D=8
M506 23626 23628 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=468970 $D=8
M507 24146 23884 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=70365 $Y=112830 $D=8
M508 23932 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=70720 $Y=160970 $D=8
M509 23931 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=70720 $Y=164845 $D=8
M510 VDD 23454 23456 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=179690 $D=8
M511 VDD 24203 24202 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=180970 $D=8
M512 VDD 24211 24210 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=323690 $D=8
M513 VDD 24219 24218 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=324970 $D=8
M514 VDD 24227 24226 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=467690 $D=8
M515 VDD 23622 23624 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=468970 $D=8
M516 23454 23456 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=179690 $D=8
M517 24203 24202 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=180970 $D=8
M518 24211 24210 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=323690 $D=8
M519 24219 24218 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=324970 $D=8
M520 24227 24226 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=467690 $D=8
M521 23622 23624 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=468970 $D=8
M522 23933 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=73815 $Y=160970 $D=8
M523 23934 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=73815 $Y=164845 $D=8
M524 24147 23883 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=74030 $Y=112830 $D=8
M525 VDD 23450 23452 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=179690 $D=8
M526 VDD 24205 24204 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=180970 $D=8
M527 VDD 24213 24212 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=323690 $D=8
M528 VDD 24221 24220 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=324970 $D=8
M529 VDD 24229 24228 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=467690 $D=8
M530 VDD 23618 23620 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=468970 $D=8
M531 23450 23452 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=179690 $D=8
M532 24205 24204 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=180970 $D=8
M533 24213 24212 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=323690 $D=8
M534 24221 24220 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=324970 $D=8
M535 24229 24228 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=467690 $D=8
M536 23618 23620 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=468970 $D=8
M537 24148 23882 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=76560 $Y=112830 $D=8
M538 23936 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=76915 $Y=160970 $D=8
M539 23935 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=76915 $Y=164845 $D=8
M540 VDD 23358 23360 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=179690 $D=8
M541 VDD 24359 24358 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=180970 $D=8
M542 VDD 24383 24382 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=323690 $D=8
M543 VDD 24407 24406 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=324970 $D=8
M544 VDD 24431 24430 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=467690 $D=8
M545 VDD 23614 23616 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=468970 $D=8
M546 23358 23360 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=179690 $D=8
M547 24359 24358 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=180970 $D=8
M548 24383 24382 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=323690 $D=8
M549 24407 24406 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=324970 $D=8
M550 24431 24430 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=467690 $D=8
M551 23614 23616 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=468970 $D=8
M552 23937 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=80005 $Y=160970 $D=8
M553 23938 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=80005 $Y=164845 $D=8
M554 24149 23881 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=80220 $Y=112830 $D=8
M555 VDD 23354 23356 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=179690 $D=8
M556 VDD 24361 24360 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=180970 $D=8
M557 VDD 24385 24384 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=323690 $D=8
M558 VDD 24409 24408 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=324970 $D=8
M559 VDD 24433 24432 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=467690 $D=8
M560 VDD 23610 23612 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=468970 $D=8
M561 23354 23356 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=179690 $D=8
M562 24361 24360 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=180970 $D=8
M563 24385 24384 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=323690 $D=8
M564 24409 24408 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=324970 $D=8
M565 24433 24432 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=467690 $D=8
M566 23610 23612 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=468970 $D=8
M567 24150 23880 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=82750 $Y=112830 $D=8
M568 23940 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=83105 $Y=160970 $D=8
M569 23939 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=83105 $Y=164845 $D=8
M570 VDD 23366 23368 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=179690 $D=8
M571 VDD 24363 24362 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=180970 $D=8
M572 VDD 24387 24386 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=323690 $D=8
M573 VDD 24411 24410 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=324970 $D=8
M574 VDD 24435 24434 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=467690 $D=8
M575 VDD 23606 23608 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=468970 $D=8
M576 23366 23368 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=179690 $D=8
M577 24363 24362 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=180970 $D=8
M578 24387 24386 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=323690 $D=8
M579 24411 24410 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=324970 $D=8
M580 24435 24434 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=467690 $D=8
M581 23606 23608 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=468970 $D=8
M582 23941 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=86200 $Y=160970 $D=8
M583 23942 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=86200 $Y=164845 $D=8
M584 24151 23879 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=86415 $Y=112830 $D=8
M585 VDD 23362 23364 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=179690 $D=8
M586 VDD 24365 24364 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=180970 $D=8
M587 VDD 24389 24388 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=323690 $D=8
M588 VDD 24413 24412 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=324970 $D=8
M589 VDD 24437 24436 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=467690 $D=8
M590 VDD 23602 23604 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=468970 $D=8
M591 23362 23364 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=179690 $D=8
M592 24365 24364 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=180970 $D=8
M593 24389 24388 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=323690 $D=8
M594 24413 24412 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=324970 $D=8
M595 24437 24436 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=467690 $D=8
M596 23602 23604 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=468970 $D=8
M597 24035 23878 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=88945 $Y=112830 $D=8
M598 1066 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=89120 $Y=160970 $D=8
M599 1067 23199 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=89120 $Y=164845 $D=8
M600 1079 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=92575 $Y=160970 $D=8
M601 1080 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=92575 $Y=164845 $D=8
M602 VDD 23662 23664 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=179690 $D=8
M603 VDD 24380 24381 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=180970 $D=8
M604 VDD 24404 24405 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=323690 $D=8
M605 VDD 24428 24429 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=324970 $D=8
M606 VDD 24452 24453 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=467690 $D=8
M607 VDD 23694 23696 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=468970 $D=8
M608 24039 23885 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=92620 $Y=112830 $D=8
M609 23662 23664 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=179690 $D=8
M610 24380 24381 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=180970 $D=8
M611 24404 24405 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=323690 $D=8
M612 24428 24429 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=324970 $D=8
M613 24452 24453 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=467690 $D=8
M614 23694 23696 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=468970 $D=8
M615 24659 23884 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=95145 $Y=112830 $D=8
M616 23997 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=95500 $Y=160970 $D=8
M617 23998 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=95500 $Y=164845 $D=8
M618 VDD 23658 23660 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=179690 $D=8
M619 VDD 24378 24379 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=180970 $D=8
M620 VDD 24402 24403 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=323690 $D=8
M621 VDD 24426 24427 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=324970 $D=8
M622 VDD 24450 24451 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=467690 $D=8
M623 VDD 23690 23692 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=468970 $D=8
M624 23658 23660 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=179690 $D=8
M625 24378 24379 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=180970 $D=8
M626 24402 24403 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=323690 $D=8
M627 24426 24427 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=324970 $D=8
M628 24450 24451 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=467690 $D=8
M629 23690 23692 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=468970 $D=8
M630 23996 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=98595 $Y=160970 $D=8
M631 23995 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=98595 $Y=164845 $D=8
M632 VDD 23654 23656 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=179690 $D=8
M633 VDD 24376 24377 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=180970 $D=8
M634 VDD 24400 24401 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=323690 $D=8
M635 VDD 24424 24425 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=324970 $D=8
M636 VDD 24448 24449 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=467690 $D=8
M637 VDD 23686 23688 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=468970 $D=8
M638 24658 23883 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=98810 $Y=112830 $D=8
M639 23654 23656 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=179690 $D=8
M640 24376 24377 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=180970 $D=8
M641 24400 24401 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=323690 $D=8
M642 24424 24425 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=324970 $D=8
M643 24448 24449 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=467690 $D=8
M644 23686 23688 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=468970 $D=8
M645 24657 23882 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=101340 $Y=112830 $D=8
M646 23993 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=101695 $Y=160970 $D=8
M647 23994 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=101695 $Y=164845 $D=8
M648 VDD 23650 23652 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=179690 $D=8
M649 VDD 24374 24375 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=180970 $D=8
M650 VDD 24398 24399 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=323690 $D=8
M651 VDD 24422 24423 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=324970 $D=8
M652 VDD 24446 24447 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=467690 $D=8
M653 VDD 23682 23684 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=468970 $D=8
M654 23650 23652 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=179690 $D=8
M655 24374 24375 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=180970 $D=8
M656 24398 24399 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=323690 $D=8
M657 24422 24423 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=324970 $D=8
M658 24446 24447 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=467690 $D=8
M659 23682 23684 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=468970 $D=8
M660 VDD 23646 23648 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=179690 $D=8
M661 VDD 24372 24373 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=180970 $D=8
M662 VDD 24396 24397 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=323690 $D=8
M663 VDD 24420 24421 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=324970 $D=8
M664 VDD 24444 24445 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=467690 $D=8
M665 VDD 23678 23680 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=468970 $D=8
M666 23992 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=104785 $Y=160970 $D=8
M667 23991 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=104785 $Y=164845 $D=8
M668 24656 23881 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=105000 $Y=112830 $D=8
M669 23646 23648 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=179690 $D=8
M670 24372 24373 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=180970 $D=8
M671 24396 24397 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=323690 $D=8
M672 24420 24421 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=324970 $D=8
M673 24444 24445 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=467690 $D=8
M674 23678 23680 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=468970 $D=8
M675 24655 23880 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=107530 $Y=112830 $D=8
M676 VDD 23642 23644 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=179690 $D=8
M677 VDD 24370 24371 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=180970 $D=8
M678 VDD 24394 24395 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=323690 $D=8
M679 VDD 24418 24419 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=324970 $D=8
M680 VDD 24442 24443 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=467690 $D=8
M681 VDD 23674 23676 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=468970 $D=8
M682 23989 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=107885 $Y=160970 $D=8
M683 23990 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=107885 $Y=164845 $D=8
M684 23642 23644 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=179690 $D=8
M685 24370 24371 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=180970 $D=8
M686 24394 24395 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=323690 $D=8
M687 24418 24419 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=324970 $D=8
M688 24442 24443 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=467690 $D=8
M689 23674 23676 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=468970 $D=8
M690 VDD 23638 23640 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=179690 $D=8
M691 VDD 24368 24369 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=180970 $D=8
M692 VDD 24392 24393 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=323690 $D=8
M693 VDD 24416 24417 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=324970 $D=8
M694 VDD 24440 24441 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=467690 $D=8
M695 VDD 23670 23672 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=468970 $D=8
M696 23988 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=110980 $Y=160970 $D=8
M697 23987 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=110980 $Y=164845 $D=8
M698 24654 23879 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=111195 $Y=112830 $D=8
M699 23638 23640 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=179690 $D=8
M700 24368 24369 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=180970 $D=8
M701 24392 24393 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=323690 $D=8
M702 24416 24417 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=324970 $D=8
M703 24440 24441 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=467690 $D=8
M704 23670 23672 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=468970 $D=8
M705 VDD 23634 23636 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=179690 $D=8
M706 VDD 24366 24367 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=180970 $D=8
M707 VDD 24390 24391 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=323690 $D=8
M708 VDD 24414 24415 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=324970 $D=8
M709 VDD 24438 24439 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=467690 $D=8
M710 VDD 23666 23668 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=468970 $D=8
M711 24653 23878 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=113725 $Y=112830 $D=8
M712 23985 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=114080 $Y=160970 $D=8
M713 23986 1078 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=114080 $Y=164845 $D=8
M714 23634 23636 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=179690 $D=8
M715 24366 24367 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=180970 $D=8
M716 24390 24391 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=323690 $D=8
M717 24414 24415 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=324970 $D=8
M718 24438 24439 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=467690 $D=8
M719 23666 23668 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=468970 $D=8
M720 VDD 23497 23498 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=179690 $D=8
M721 VDD 24674 24675 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=180970 $D=8
M722 VDD 24676 24677 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=215690 $D=8
M723 VDD 24678 24679 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=216970 $D=8
M724 VDD 24680 24681 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=251690 $D=8
M725 VDD 24682 24683 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=252970 $D=8
M726 VDD 24684 24685 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=287690 $D=8
M727 VDD 24686 24687 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=288970 $D=8
M728 VDD 24688 24689 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=323690 $D=8
M729 VDD 24690 24691 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=324970 $D=8
M730 VDD 24692 24693 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=359690 $D=8
M731 VDD 24694 24695 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=360970 $D=8
M732 VDD 24696 24697 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=395690 $D=8
M733 VDD 24698 24699 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=396970 $D=8
M734 VDD 24700 24701 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=431690 $D=8
M735 VDD 24702 24703 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=432970 $D=8
M736 VDD 24704 24705 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=467690 $D=8
M737 VDD 23499 23500 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=468970 $D=8
M738 VDD VSS VDD VDD pfet_05v0 L=2.365e-06 W=8.19e-05 AD=0 AS=6.1309e-11 PD=0 PS=0.000217698 NRD=0 NRS=11.8457 m=1 nf=36 $X=10835 $Y=171065 $D=8
M739 23497 23498 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=179690 $D=8
M740 24674 24675 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=180970 $D=8
M741 24676 24677 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=215690 $D=8
M742 24678 24679 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=216970 $D=8
M743 24680 24681 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=251690 $D=8
M744 24682 24683 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=252970 $D=8
M745 24684 24685 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=287690 $D=8
M746 24686 24687 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=288970 $D=8
M747 24688 24689 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=323690 $D=8
M748 24690 24691 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=324970 $D=8
M749 24692 24693 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=359690 $D=8
M750 24694 24695 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=360970 $D=8
M751 24696 24697 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=395690 $D=8
M752 24698 24699 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=396970 $D=8
M753 24700 24701 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=431690 $D=8
M754 24702 24703 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=432970 $D=8
M755 24704 24705 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=467690 $D=8
M756 23499 23500 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=468970 $D=8
M757 VDD VSS VDD VDD pfet_05v0 L=3.94e-06 W=0.000357175 AD=0 AS=2.0381e-10 PD=0 PS=0.00079952 NRD=0 NRS=6.74977 m=1 nf=65 $X=146370 $Y=180915 $D=8
M758 VDD 24106 23202 VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=156680 $Y=180895 $D=8
M759 23209 24108 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=213535 $D=8
M760 VDD 24110 23210 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=216895 $D=8
M761 23217 24112 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=249535 $D=8
M762 VDD 24114 23218 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=252895 $D=8
M763 23225 24116 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=285535 $D=8
M764 VDD 24118 23226 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=288895 $D=8
M765 23233 24120 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=321535 $D=8
M766 VDD 24122 23234 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=324895 $D=8
M767 23241 24124 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=357535 $D=8
M768 VDD 24126 23242 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=360895 $D=8
M769 23249 24128 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=393535 $D=8
M770 VDD 24130 23250 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=396895 $D=8
M771 23257 24132 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=429535 $D=8
M772 VDD 24134 23258 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=432895 $D=8
M773 23265 24136 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=156680 $Y=465535 $D=8
M774 24043 1040 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=180895 $D=8
M775 VDD 1044 24043 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=182015 $D=8
M776 24043 1052 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=183135 $D=8
M777 VDD 1045 24045 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=213535 $D=8
M778 24045 1044 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=214655 $D=8
M779 VDD 1040 24045 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=215775 $D=8
M780 24047 1040 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=216895 $D=8
M781 VDD 1043 24047 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=218015 $D=8
M782 24047 1052 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=219135 $D=8
M783 VDD 1045 24049 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=249535 $D=8
M784 24049 1043 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=250655 $D=8
M785 VDD 1040 24049 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=251775 $D=8
M786 24051 1040 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=252895 $D=8
M787 VDD 1042 24051 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=254015 $D=8
M788 24051 1052 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=255135 $D=8
M789 VDD 1045 24053 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=285535 $D=8
M790 24053 1042 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=286655 $D=8
M791 VDD 1040 24053 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=287775 $D=8
M792 24055 1040 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=288895 $D=8
M793 VDD 1041 24055 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=290015 $D=8
M794 24055 1052 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=291135 $D=8
M795 VDD 1045 24057 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=321535 $D=8
M796 24057 1041 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=322655 $D=8
M797 VDD 1040 24057 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=323775 $D=8
M798 24059 1038 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=324895 $D=8
M799 VDD 1044 24059 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=326015 $D=8
M800 24059 1052 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=327135 $D=8
M801 VDD 1045 24061 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=357535 $D=8
M802 24061 1044 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=358655 $D=8
M803 VDD 1038 24061 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=359775 $D=8
M804 24063 1038 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=360895 $D=8
M805 VDD 1043 24063 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=362015 $D=8
M806 24063 1052 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=363135 $D=8
M807 VDD 1045 24065 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=393535 $D=8
M808 24065 1043 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=394655 $D=8
M809 VDD 1038 24065 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=395775 $D=8
M810 24067 1038 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=396895 $D=8
M811 VDD 1042 24067 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=398015 $D=8
M812 24067 1052 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=399135 $D=8
M813 VDD 1045 24069 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=429535 $D=8
M814 24069 1042 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=430655 $D=8
M815 VDD 1038 24069 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=431775 $D=8
M816 24071 1038 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=432895 $D=8
M817 VDD 1041 24071 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=434015 $D=8
M818 24071 1052 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=435135 $D=8
M819 VDD 1045 24073 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=465535 $D=8
M820 24073 1041 VDD VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=466655 $D=8
M821 VDD 1038 24073 VDD pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=467775 $D=8
M822 24033 1 VDD VDD pfet_05v0 L=5.95e-07 W=2.28e-06 AD=5.985e-13 AS=1.3566e-12 PD=2.805e-06 PS=5.75e-06 NRD=0.115132 NRS=0.260965 m=1 nf=1 $X=233770 $Y=57780 $D=8
M823 617 1000 VDD VDD pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=233770 $Y=63100 $D=8
M824 1000 CLK 24033 VDD pfet_05v0 L=5.95e-07 W=2.28e-06 AD=1.3566e-12 AS=5.985e-13 PD=5.75e-06 PS=2.805e-06 NRD=0.260965 NRS=0.115132 m=1 nf=1 $X=234890 $Y=57780 $D=8
M825 616 619 VDD VDD pfet_05v0 L=6e-07 W=1.134e-05 AD=2.9484e-12 AS=4.9896e-12 PD=1.238e-05 PS=2.444e-05 NRD=0.0917108 NRS=0.155203 m=1 nf=2 $X=242235 $Y=57810 $D=8
M826 281 1006 VDD VDD pfet_05v0 L=1e-06 W=9e-07 AD=3.96e-13 AS=3.96e-13 PD=2.68e-06 PS=2.68e-06 NRD=0.488889 NRS=0.488889 m=1 nf=1 $X=243265 $Y=42525 $D=8
M827 CEN 617 619 VDD pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=245925 $Y=59010 $D=8
M828 618 1000 619 VDD pfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=245925 $Y=64875 $D=8
M829 317 281 VDD VDD pfet_05v0 L=6e-07 W=1.89e-06 AD=8.316e-13 AS=8.316e-13 PD=4.66e-06 PS=4.66e-06 NRD=0.232804 NRS=0.232804 m=1 nf=1 $X=246495 $Y=41535 $D=8
M830 354 317 VDD VDD pfet_05v0 L=6e-07 W=7.54e-06 AD=1.9604e-12 AS=3.3176e-12 PD=8.58e-06 PS=1.684e-05 NRD=0.137931 NRS=0.233422 m=1 nf=2 $X=249065 $Y=39655 $D=8
M831 250 468 VDD VDD pfet_05v0 L=6e-07 W=0.0001248 AD=3.2448e-11 AS=3.69283e-11 PD=0.00013 PS=0.000130718 NRD=0.208333 NRS=0.237099 m=1 nf=10 $X=240535 $Y=94430 $D=8
M832 445 354 VDD VDD pfet_05v0 L=6e-07 W=1.95e-05 AD=5.07e-12 AS=8.58e-12 PD=2.002e-05 PS=3.988e-05 NRD=0.0133333 NRS=0.0225641 m=1 nf=1 $X=256125 $Y=53590 $D=8
M833 VDD CLK 445 VDD pfet_05v0 L=6e-07 W=1.95e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=257245 $Y=53590 $D=8
M834 445 616 VDD VDD pfet_05v0 L=6e-07 W=1.95e-05 AD=8.58e-12 AS=5.07e-12 PD=3.988e-05 PS=2.002e-05 NRD=0.0225641 NRS=0.0133333 m=1 nf=1 $X=258365 $Y=53590 $D=8
M835 VDD 495 468 VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=9.9792e-12 PD=2.32e-05 PS=4.624e-05 NRD=0.0114638 NRS=0.0194004 m=1 nf=1 $X=262120 $Y=50420 $D=8
M836 468 445 VDD VDD pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.64e-05 PS=4.64e-05 NRD=0.0229277 NRS=0.0229277 m=1 nf=2 $X=263240 $Y=50420 $D=8
M837 468 495 VDD VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=9.9792e-12 AS=5.8968e-12 PD=4.624e-05 PS=2.32e-05 NRD=0.0194004 NRS=0.0114638 m=1 nf=1 $X=265480 $Y=50420 $D=8
M838 VDD 24107 23266 VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=258945 $Y=180895 $D=8
M839 23273 24109 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=213535 $D=8
M840 VDD 24111 23274 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=216895 $D=8
M841 23281 24113 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=249535 $D=8
M842 VDD 24115 23282 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=252895 $D=8
M843 23289 24117 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=285535 $D=8
M844 VDD 24119 23290 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=288895 $D=8
M845 23297 24121 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=321535 $D=8
M846 VDD 24123 23298 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=324895 $D=8
M847 23305 24125 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=357535 $D=8
M848 VDD 24127 23306 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=360895 $D=8
M849 23313 24129 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=393535 $D=8
M850 VDD 24131 23314 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=396895 $D=8
M851 23321 24133 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=429535 $D=8
M852 VDD 24135 23322 VDD pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=432895 $D=8
M853 23329 24137 VDD VDD pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=258945 $Y=465535 $D=8
M854 VDD 468 495 VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=9.9792e-12 PD=2.32e-05 PS=4.624e-05 NRD=0.0114638 NRS=0.0194004 m=1 nf=1 $X=268545 $Y=50420 $D=8
M855 495 607 VDD VDD pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.64e-05 PS=4.64e-05 NRD=0.0229277 NRS=0.0229277 m=1 nf=2 $X=269665 $Y=50420 $D=8
M856 495 468 VDD VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=9.9792e-12 AS=5.8968e-12 PD=4.624e-05 PS=2.32e-05 NRD=0.0194004 NRS=0.0114638 m=1 nf=1 $X=271905 $Y=50420 $D=8
M857 1 250 VDD VDD pfet_05v0 L=6e-07 W=0.0003674 AD=9.5524e-11 AS=1.02119e-10 PD=0.0003778 PS=0.000378518 NRD=0.28307 NRS=0.302613 m=1 nf=20 $X=253180 $Y=88540 $D=8
M858 VDD VSS VDD VDD pfet_05v0 L=3.94e-06 W=0.000357175 AD=0 AS=2.0381e-10 PD=0 PS=0.00079952 NRD=0 NRS=6.74977 m=1 nf=65 $X=273750 $Y=180915 $D=8
M859 VDD 23501 23502 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=179690 $D=8
M860 VDD 24754 24755 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=180970 $D=8
M861 VDD 24756 24757 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=215690 $D=8
M862 VDD 24774 24775 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=216970 $D=8
M863 VDD 24776 24777 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=251690 $D=8
M864 VDD 24794 24795 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=252970 $D=8
M865 VDD 24796 24797 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=287690 $D=8
M866 VDD 24814 24815 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=288970 $D=8
M867 VDD 24816 24817 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=323690 $D=8
M868 VDD 24834 24835 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=324970 $D=8
M869 VDD 24836 24837 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=359690 $D=8
M870 VDD 24854 24855 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=360970 $D=8
M871 VDD 24856 24857 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=395690 $D=8
M872 VDD 24874 24875 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=396970 $D=8
M873 VDD 24876 24877 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=431690 $D=8
M874 VDD 24894 24895 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=432970 $D=8
M875 VDD 24896 24897 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=467690 $D=8
M876 VDD 23503 23504 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=468970 $D=8
M877 23501 23502 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=179690 $D=8
M878 24754 24755 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=180970 $D=8
M879 24756 24757 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=215690 $D=8
M880 24774 24775 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=216970 $D=8
M881 24776 24777 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=251690 $D=8
M882 24794 24795 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=252970 $D=8
M883 24796 24797 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=287690 $D=8
M884 24814 24815 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=288970 $D=8
M885 24816 24817 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=323690 $D=8
M886 24834 24835 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=324970 $D=8
M887 24836 24837 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=359690 $D=8
M888 24854 24855 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=360970 $D=8
M889 24856 24857 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=395690 $D=8
M890 24874 24875 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=396970 $D=8
M891 24876 24877 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=431690 $D=8
M892 24894 24895 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=432970 $D=8
M893 24896 24897 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=467690 $D=8
M894 23503 23504 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=468970 $D=8
M895 VDD 23478 23480 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=179690 $D=8
M896 VDD 24739 24738 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=180970 $D=8
M897 VDD 24747 24746 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=215690 $D=8
M898 VDD 24759 24758 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=216970 $D=8
M899 VDD 24767 24766 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=251690 $D=8
M900 VDD 24779 24778 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=252970 $D=8
M901 VDD 24787 24786 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=287690 $D=8
M902 VDD 24799 24798 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=288970 $D=8
M903 VDD 24807 24806 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=323690 $D=8
M904 VDD 24819 24818 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=324970 $D=8
M905 VDD 24827 24826 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=359690 $D=8
M906 VDD 24839 24838 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=360970 $D=8
M907 VDD 24847 24846 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=395690 $D=8
M908 VDD 24859 24858 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=396970 $D=8
M909 VDD 24867 24866 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=431690 $D=8
M910 VDD 24879 24878 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=432970 $D=8
M911 VDD 24887 24886 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=467690 $D=8
M912 VDD 23414 23416 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=468970 $D=8
M913 23478 23480 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=179690 $D=8
M914 24739 24738 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=180970 $D=8
M915 24747 24746 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=215690 $D=8
M916 24759 24758 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=216970 $D=8
M917 24767 24766 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=251690 $D=8
M918 24779 24778 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=252970 $D=8
M919 24787 24786 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=287690 $D=8
M920 24799 24798 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=288970 $D=8
M921 24807 24806 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=323690 $D=8
M922 24819 24818 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=324970 $D=8
M923 24827 24826 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=359690 $D=8
M924 24839 24838 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=360970 $D=8
M925 24847 24846 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=395690 $D=8
M926 24859 24858 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=396970 $D=8
M927 24867 24866 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=431690 $D=8
M928 24879 24878 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=432970 $D=8
M929 24887 24886 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=467690 $D=8
M930 23414 23416 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=468970 $D=8
M931 23943 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=311500 $Y=160970 $D=8
M932 23944 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=311500 $Y=164845 $D=8
M933 24152 23886 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=311715 $Y=112830 $D=8
M934 VDD 23474 23476 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=179690 $D=8
M935 VDD 24741 24740 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=180970 $D=8
M936 VDD 24749 24748 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=215690 $D=8
M937 VDD 24761 24760 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=216970 $D=8
M938 VDD 24769 24768 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=251690 $D=8
M939 VDD 24781 24780 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=252970 $D=8
M940 VDD 24789 24788 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=287690 $D=8
M941 VDD 24801 24800 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=288970 $D=8
M942 VDD 24809 24808 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=323690 $D=8
M943 VDD 24821 24820 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=324970 $D=8
M944 VDD 24829 24828 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=359690 $D=8
M945 VDD 24841 24840 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=360970 $D=8
M946 VDD 24849 24848 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=395690 $D=8
M947 VDD 24861 24860 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=396970 $D=8
M948 VDD 24869 24868 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=431690 $D=8
M949 VDD 24881 24880 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=432970 $D=8
M950 VDD 24889 24888 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=467690 $D=8
M951 VDD 23410 23412 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=468970 $D=8
M952 23474 23476 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=179690 $D=8
M953 24741 24740 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=180970 $D=8
M954 24749 24748 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=215690 $D=8
M955 24761 24760 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=216970 $D=8
M956 24769 24768 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=251690 $D=8
M957 24781 24780 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=252970 $D=8
M958 24789 24788 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=287690 $D=8
M959 24801 24800 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=288970 $D=8
M960 24809 24808 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=323690 $D=8
M961 24821 24820 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=324970 $D=8
M962 24829 24828 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=359690 $D=8
M963 24841 24840 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=360970 $D=8
M964 24849 24848 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=395690 $D=8
M965 24861 24860 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=396970 $D=8
M966 24869 24868 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=431690 $D=8
M967 24881 24880 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=432970 $D=8
M968 24889 24888 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=467690 $D=8
M969 23410 23412 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=468970 $D=8
M970 24153 23887 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=314245 $Y=112830 $D=8
M971 23946 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=314600 $Y=160970 $D=8
M972 23945 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=314600 $Y=164845 $D=8
M973 VDD 23470 23472 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=179690 $D=8
M974 VDD 24743 24742 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=180970 $D=8
M975 VDD 24751 24750 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=215690 $D=8
M976 VDD 24763 24762 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=216970 $D=8
M977 VDD 24771 24770 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=251690 $D=8
M978 VDD 24783 24782 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=252970 $D=8
M979 VDD 24791 24790 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=287690 $D=8
M980 VDD 24803 24802 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=288970 $D=8
M981 VDD 24811 24810 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=323690 $D=8
M982 VDD 24823 24822 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=324970 $D=8
M983 VDD 24831 24830 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=359690 $D=8
M984 VDD 24843 24842 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=360970 $D=8
M985 VDD 24851 24850 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=395690 $D=8
M986 VDD 24863 24862 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=396970 $D=8
M987 VDD 24871 24870 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=431690 $D=8
M988 VDD 24883 24882 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=432970 $D=8
M989 VDD 24891 24890 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=467690 $D=8
M990 VDD 23406 23408 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=468970 $D=8
M991 23470 23472 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=179690 $D=8
M992 24743 24742 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=180970 $D=8
M993 24751 24750 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=215690 $D=8
M994 24763 24762 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=216970 $D=8
M995 24771 24770 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=251690 $D=8
M996 24783 24782 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=252970 $D=8
M997 24791 24790 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=287690 $D=8
M998 24803 24802 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=288970 $D=8
M999 24811 24810 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=323690 $D=8
M1000 24823 24822 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=324970 $D=8
M1001 24831 24830 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=359690 $D=8
M1002 24843 24842 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=360970 $D=8
M1003 24851 24850 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=395690 $D=8
M1004 24863 24862 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=396970 $D=8
M1005 24871 24870 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=431690 $D=8
M1006 24883 24882 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=432970 $D=8
M1007 24891 24890 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=467690 $D=8
M1008 23406 23408 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=468970 $D=8
M1009 23947 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=317695 $Y=160970 $D=8
M1010 23948 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=317695 $Y=164845 $D=8
M1011 24154 23888 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=317910 $Y=112830 $D=8
M1012 VDD 23466 23468 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=179690 $D=8
M1013 VDD 24745 24744 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=180970 $D=8
M1014 VDD 24753 24752 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=215690 $D=8
M1015 VDD 24765 24764 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=216970 $D=8
M1016 VDD 24773 24772 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=251690 $D=8
M1017 VDD 24785 24784 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=252970 $D=8
M1018 VDD 24793 24792 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=287690 $D=8
M1019 VDD 24805 24804 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=288970 $D=8
M1020 VDD 24813 24812 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=323690 $D=8
M1021 VDD 24825 24824 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=324970 $D=8
M1022 VDD 24833 24832 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=359690 $D=8
M1023 VDD 24845 24844 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=360970 $D=8
M1024 VDD 24853 24852 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=395690 $D=8
M1025 VDD 24865 24864 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=396970 $D=8
M1026 VDD 24873 24872 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=431690 $D=8
M1027 VDD 24885 24884 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=432970 $D=8
M1028 VDD 24893 24892 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=467690 $D=8
M1029 VDD 23402 23404 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=468970 $D=8
M1030 23466 23468 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=179690 $D=8
M1031 24745 24744 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=180970 $D=8
M1032 24753 24752 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=215690 $D=8
M1033 24765 24764 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=216970 $D=8
M1034 24773 24772 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=251690 $D=8
M1035 24785 24784 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=252970 $D=8
M1036 24793 24792 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=287690 $D=8
M1037 24805 24804 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=288970 $D=8
M1038 24813 24812 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=323690 $D=8
M1039 24825 24824 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=324970 $D=8
M1040 24833 24832 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=359690 $D=8
M1041 24845 24844 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=360970 $D=8
M1042 24853 24852 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=395690 $D=8
M1043 24865 24864 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=396970 $D=8
M1044 24873 24872 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=431690 $D=8
M1045 24885 24884 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=432970 $D=8
M1046 24893 24892 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=467690 $D=8
M1047 23402 23404 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=468970 $D=8
M1048 24155 23889 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=320440 $Y=112830 $D=8
M1049 23950 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=320795 $Y=160970 $D=8
M1050 23949 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=320795 $Y=164845 $D=8
M1051 VDD 23374 23376 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=179690 $D=8
M1052 VDD 24455 24454 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=180970 $D=8
M1053 VDD 24479 24478 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=323690 $D=8
M1054 VDD 24503 24502 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=324970 $D=8
M1055 VDD 24527 24526 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=467690 $D=8
M1056 VDD 23430 23432 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=468970 $D=8
M1057 23374 23376 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=179690 $D=8
M1058 24455 24454 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=180970 $D=8
M1059 24479 24478 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=323690 $D=8
M1060 24503 24502 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=324970 $D=8
M1061 24527 24526 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=467690 $D=8
M1062 23430 23432 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=468970 $D=8
M1063 23951 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=323885 $Y=160970 $D=8
M1064 23952 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=323885 $Y=164845 $D=8
M1065 24156 23890 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=324100 $Y=112830 $D=8
M1066 VDD 23370 23372 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=179690 $D=8
M1067 VDD 24457 24456 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=180970 $D=8
M1068 VDD 24481 24480 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=323690 $D=8
M1069 VDD 24505 24504 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=324970 $D=8
M1070 VDD 24529 24528 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=467690 $D=8
M1071 VDD 23426 23428 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=468970 $D=8
M1072 23370 23372 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=179690 $D=8
M1073 24457 24456 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=180970 $D=8
M1074 24481 24480 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=323690 $D=8
M1075 24505 24504 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=324970 $D=8
M1076 24529 24528 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=467690 $D=8
M1077 23426 23428 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=468970 $D=8
M1078 24157 23891 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=326630 $Y=112830 $D=8
M1079 23954 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=326985 $Y=160970 $D=8
M1080 23953 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=326985 $Y=164845 $D=8
M1081 VDD 23382 23384 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=179690 $D=8
M1082 VDD 24459 24458 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=180970 $D=8
M1083 VDD 24483 24482 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=323690 $D=8
M1084 VDD 24507 24506 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=324970 $D=8
M1085 VDD 24531 24530 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=467690 $D=8
M1086 VDD 23422 23424 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=468970 $D=8
M1087 23382 23384 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=179690 $D=8
M1088 24459 24458 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=180970 $D=8
M1089 24483 24482 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=323690 $D=8
M1090 24507 24506 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=324970 $D=8
M1091 24531 24530 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=467690 $D=8
M1092 23422 23424 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=468970 $D=8
M1093 23955 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=330080 $Y=160970 $D=8
M1094 23956 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=330080 $Y=164845 $D=8
M1095 24158 23892 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=330295 $Y=112830 $D=8
M1096 VDD 23378 23380 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=179690 $D=8
M1097 VDD 24461 24460 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=180970 $D=8
M1098 VDD 24485 24484 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=323690 $D=8
M1099 VDD 24509 24508 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=324970 $D=8
M1100 VDD 24533 24532 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=467690 $D=8
M1101 VDD 23418 23420 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=468970 $D=8
M1102 23378 23380 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=179690 $D=8
M1103 24461 24460 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=180970 $D=8
M1104 24485 24484 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=323690 $D=8
M1105 24509 24508 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=324970 $D=8
M1106 24533 24532 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=467690 $D=8
M1107 23418 23420 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=468970 $D=8
M1108 24036 23893 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=332825 $Y=112830 $D=8
M1109 1069 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=333000 $Y=160970 $D=8
M1110 1070 23200 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=333000 $Y=164845 $D=8
M1111 1083 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=336455 $Y=160970 $D=8
M1112 1084 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=336455 $Y=164845 $D=8
M1113 VDD 23726 23728 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=179690 $D=8
M1114 VDD 24476 24477 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=180970 $D=8
M1115 VDD 24500 24501 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=323690 $D=8
M1116 VDD 24524 24525 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=324970 $D=8
M1117 VDD 24548 24549 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=467690 $D=8
M1118 VDD 23758 23760 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=468970 $D=8
M1119 24040 23886 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=336500 $Y=112830 $D=8
M1120 23726 23728 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=179690 $D=8
M1121 24476 24477 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=180970 $D=8
M1122 24500 24501 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=323690 $D=8
M1123 24524 24525 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=324970 $D=8
M1124 24548 24549 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=467690 $D=8
M1125 23758 23760 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=468970 $D=8
M1126 24666 23887 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=339025 $Y=112830 $D=8
M1127 24011 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=339380 $Y=160970 $D=8
M1128 24012 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=339380 $Y=164845 $D=8
M1129 VDD 23722 23724 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=179690 $D=8
M1130 VDD 24474 24475 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=180970 $D=8
M1131 VDD 24498 24499 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=323690 $D=8
M1132 VDD 24522 24523 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=324970 $D=8
M1133 VDD 24546 24547 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=467690 $D=8
M1134 VDD 23754 23756 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=468970 $D=8
M1135 23722 23724 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=179690 $D=8
M1136 24474 24475 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=180970 $D=8
M1137 24498 24499 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=323690 $D=8
M1138 24522 24523 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=324970 $D=8
M1139 24546 24547 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=467690 $D=8
M1140 23754 23756 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=468970 $D=8
M1141 24010 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=342475 $Y=160970 $D=8
M1142 24009 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=342475 $Y=164845 $D=8
M1143 VDD 23718 23720 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=179690 $D=8
M1144 VDD 24472 24473 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=180970 $D=8
M1145 VDD 24496 24497 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=323690 $D=8
M1146 VDD 24520 24521 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=324970 $D=8
M1147 VDD 24544 24545 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=467690 $D=8
M1148 VDD 23750 23752 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=468970 $D=8
M1149 24665 23888 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=342690 $Y=112830 $D=8
M1150 23718 23720 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=179690 $D=8
M1151 24472 24473 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=180970 $D=8
M1152 24496 24497 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=323690 $D=8
M1153 24520 24521 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=324970 $D=8
M1154 24544 24545 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=467690 $D=8
M1155 23750 23752 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=468970 $D=8
M1156 24664 23889 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=345220 $Y=112830 $D=8
M1157 24007 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=345575 $Y=160970 $D=8
M1158 24008 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=345575 $Y=164845 $D=8
M1159 VDD 23714 23716 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=179690 $D=8
M1160 VDD 24470 24471 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=180970 $D=8
M1161 VDD 24494 24495 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=323690 $D=8
M1162 VDD 24518 24519 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=324970 $D=8
M1163 VDD 24542 24543 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=467690 $D=8
M1164 VDD 23746 23748 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=468970 $D=8
M1165 23714 23716 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=179690 $D=8
M1166 24470 24471 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=180970 $D=8
M1167 24494 24495 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=323690 $D=8
M1168 24518 24519 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=324970 $D=8
M1169 24542 24543 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=467690 $D=8
M1170 23746 23748 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=468970 $D=8
M1171 VDD 23710 23712 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=179690 $D=8
M1172 VDD 24468 24469 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=180970 $D=8
M1173 VDD 24492 24493 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=323690 $D=8
M1174 VDD 24516 24517 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=324970 $D=8
M1175 VDD 24540 24541 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=467690 $D=8
M1176 VDD 23742 23744 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=468970 $D=8
M1177 24006 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=348665 $Y=160970 $D=8
M1178 24005 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=348665 $Y=164845 $D=8
M1179 24663 23890 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=348880 $Y=112830 $D=8
M1180 23710 23712 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=179690 $D=8
M1181 24468 24469 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=180970 $D=8
M1182 24492 24493 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=323690 $D=8
M1183 24516 24517 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=324970 $D=8
M1184 24540 24541 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=467690 $D=8
M1185 23742 23744 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=468970 $D=8
M1186 24662 23891 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=351410 $Y=112830 $D=8
M1187 VDD 23706 23708 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=179690 $D=8
M1188 VDD 24466 24467 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=180970 $D=8
M1189 VDD 24490 24491 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=323690 $D=8
M1190 VDD 24514 24515 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=324970 $D=8
M1191 VDD 24538 24539 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=467690 $D=8
M1192 VDD 23738 23740 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=468970 $D=8
M1193 24003 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=351765 $Y=160970 $D=8
M1194 24004 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=351765 $Y=164845 $D=8
M1195 23706 23708 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=179690 $D=8
M1196 24466 24467 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=180970 $D=8
M1197 24490 24491 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=323690 $D=8
M1198 24514 24515 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=324970 $D=8
M1199 24538 24539 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=467690 $D=8
M1200 23738 23740 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=468970 $D=8
M1201 VDD 23702 23704 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=179690 $D=8
M1202 VDD 24464 24465 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=180970 $D=8
M1203 VDD 24488 24489 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=323690 $D=8
M1204 VDD 24512 24513 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=324970 $D=8
M1205 VDD 24536 24537 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=467690 $D=8
M1206 VDD 23734 23736 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=468970 $D=8
M1207 24002 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=354860 $Y=160970 $D=8
M1208 24001 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=354860 $Y=164845 $D=8
M1209 24661 23892 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=355075 $Y=112830 $D=8
M1210 23702 23704 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=179690 $D=8
M1211 24464 24465 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=180970 $D=8
M1212 24488 24489 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=323690 $D=8
M1213 24512 24513 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=324970 $D=8
M1214 24536 24537 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=467690 $D=8
M1215 23734 23736 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=468970 $D=8
M1216 VDD 23698 23700 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=179690 $D=8
M1217 VDD 24462 24463 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=180970 $D=8
M1218 VDD 24486 24487 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=323690 $D=8
M1219 VDD 24510 24511 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=324970 $D=8
M1220 VDD 24534 24535 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=467690 $D=8
M1221 VDD 23730 23732 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=468970 $D=8
M1222 24660 23893 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=357605 $Y=112830 $D=8
M1223 23999 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=357960 $Y=160970 $D=8
M1224 24000 1081 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=357960 $Y=164845 $D=8
M1225 23698 23700 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=179690 $D=8
M1226 24462 24463 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=180970 $D=8
M1227 24486 24487 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=323690 $D=8
M1228 24510 24511 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=324970 $D=8
M1229 24534 24535 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=467690 $D=8
M1230 23730 23732 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=468970 $D=8
M1231 VDD 23494 23496 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=179690 $D=8
M1232 VDD 24231 24230 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=180970 $D=8
M1233 VDD 24239 24238 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=323690 $D=8
M1234 VDD 24247 24246 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=324970 $D=8
M1235 VDD 24255 24254 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=467690 $D=8
M1236 VDD 23790 23792 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=468970 $D=8
M1237 23494 23496 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=179690 $D=8
M1238 24231 24230 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=180970 $D=8
M1239 24239 24238 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=323690 $D=8
M1240 24247 24246 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=324970 $D=8
M1241 24255 24254 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=467690 $D=8
M1242 23790 23792 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=468970 $D=8
M1243 23957 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=365500 $Y=160970 $D=8
M1244 23958 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=365500 $Y=164845 $D=8
M1245 24159 23886 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=365715 $Y=112830 $D=8
M1246 VDD 23490 23492 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=179690 $D=8
M1247 VDD 24233 24232 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=180970 $D=8
M1248 VDD 24241 24240 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=323690 $D=8
M1249 VDD 24249 24248 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=324970 $D=8
M1250 VDD 24257 24256 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=467690 $D=8
M1251 VDD 23786 23788 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=468970 $D=8
M1252 23490 23492 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=179690 $D=8
M1253 24233 24232 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=180970 $D=8
M1254 24241 24240 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=323690 $D=8
M1255 24249 24248 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=324970 $D=8
M1256 24257 24256 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=467690 $D=8
M1257 23786 23788 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=468970 $D=8
M1258 24160 23887 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=368245 $Y=112830 $D=8
M1259 23960 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=368600 $Y=160970 $D=8
M1260 23959 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=368600 $Y=164845 $D=8
M1261 VDD 23486 23488 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=179690 $D=8
M1262 VDD 24235 24234 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=180970 $D=8
M1263 VDD 24243 24242 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=323690 $D=8
M1264 VDD 24251 24250 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=324970 $D=8
M1265 VDD 24259 24258 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=467690 $D=8
M1266 VDD 23782 23784 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=468970 $D=8
M1267 23486 23488 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=179690 $D=8
M1268 24235 24234 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=180970 $D=8
M1269 24243 24242 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=323690 $D=8
M1270 24251 24250 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=324970 $D=8
M1271 24259 24258 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=467690 $D=8
M1272 23782 23784 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=468970 $D=8
M1273 23961 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=371695 $Y=160970 $D=8
M1274 23962 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=371695 $Y=164845 $D=8
M1275 24161 23888 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=371910 $Y=112830 $D=8
M1276 VDD 23482 23484 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=179690 $D=8
M1277 VDD 24237 24236 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=180970 $D=8
M1278 VDD 24245 24244 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=323690 $D=8
M1279 VDD 24253 24252 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=324970 $D=8
M1280 VDD 24261 24260 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=467690 $D=8
M1281 VDD 23778 23780 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=468970 $D=8
M1282 23482 23484 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=179690 $D=8
M1283 24237 24236 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=180970 $D=8
M1284 24245 24244 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=323690 $D=8
M1285 24253 24252 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=324970 $D=8
M1286 24261 24260 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=467690 $D=8
M1287 23778 23780 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=468970 $D=8
M1288 24162 23889 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=374440 $Y=112830 $D=8
M1289 23964 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=374795 $Y=160970 $D=8
M1290 23963 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=374795 $Y=164845 $D=8
M1291 VDD 23390 23392 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=179690 $D=8
M1292 VDD 24551 24550 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=180970 $D=8
M1293 VDD 24575 24574 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=323690 $D=8
M1294 VDD 24599 24598 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=324970 $D=8
M1295 VDD 24623 24622 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=467690 $D=8
M1296 VDD 23774 23776 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=468970 $D=8
M1297 23390 23392 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=179690 $D=8
M1298 24551 24550 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=180970 $D=8
M1299 24575 24574 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=323690 $D=8
M1300 24599 24598 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=324970 $D=8
M1301 24623 24622 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=467690 $D=8
M1302 23774 23776 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=468970 $D=8
M1303 23965 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=377885 $Y=160970 $D=8
M1304 23966 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=377885 $Y=164845 $D=8
M1305 24163 23890 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=378100 $Y=112830 $D=8
M1306 VDD 23386 23388 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=179690 $D=8
M1307 VDD 24553 24552 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=180970 $D=8
M1308 VDD 24577 24576 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=323690 $D=8
M1309 VDD 24601 24600 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=324970 $D=8
M1310 VDD 24625 24624 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=467690 $D=8
M1311 VDD 23770 23772 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=468970 $D=8
M1312 23386 23388 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=179690 $D=8
M1313 24553 24552 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=180970 $D=8
M1314 24577 24576 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=323690 $D=8
M1315 24601 24600 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=324970 $D=8
M1316 24625 24624 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=467690 $D=8
M1317 23770 23772 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=468970 $D=8
M1318 24164 23891 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=380630 $Y=112830 $D=8
M1319 23968 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=380985 $Y=160970 $D=8
M1320 23967 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=380985 $Y=164845 $D=8
M1321 VDD 23398 23400 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=179690 $D=8
M1322 VDD 24555 24554 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=180970 $D=8
M1323 VDD 24579 24578 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=323690 $D=8
M1324 VDD 24603 24602 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=324970 $D=8
M1325 VDD 24627 24626 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=467690 $D=8
M1326 VDD 23766 23768 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=468970 $D=8
M1327 23398 23400 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=179690 $D=8
M1328 24555 24554 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=180970 $D=8
M1329 24579 24578 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=323690 $D=8
M1330 24603 24602 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=324970 $D=8
M1331 24627 24626 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=467690 $D=8
M1332 23766 23768 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=468970 $D=8
M1333 23969 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=384080 $Y=160970 $D=8
M1334 23970 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=384080 $Y=164845 $D=8
M1335 24165 23892 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=384295 $Y=112830 $D=8
M1336 VDD 23394 23396 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=179690 $D=8
M1337 VDD 24557 24556 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=180970 $D=8
M1338 VDD 24581 24580 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=323690 $D=8
M1339 VDD 24605 24604 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=324970 $D=8
M1340 VDD 24629 24628 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=467690 $D=8
M1341 VDD 23762 23764 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=468970 $D=8
M1342 23394 23396 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=179690 $D=8
M1343 24557 24556 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=180970 $D=8
M1344 24581 24580 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=323690 $D=8
M1345 24605 24604 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=324970 $D=8
M1346 24629 24628 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=467690 $D=8
M1347 23762 23764 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=468970 $D=8
M1348 24037 23893 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=386825 $Y=112830 $D=8
M1349 1072 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=387000 $Y=160970 $D=8
M1350 1073 23201 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=387000 $Y=164845 $D=8
M1351 1086 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=390455 $Y=160970 $D=8
M1352 1087 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=390455 $Y=164845 $D=8
M1353 VDD 23822 23824 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=179690 $D=8
M1354 VDD 24572 24573 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=180970 $D=8
M1355 VDD 24596 24597 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=323690 $D=8
M1356 VDD 24620 24621 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=324970 $D=8
M1357 VDD 24644 24645 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=467690 $D=8
M1358 VDD 23854 23856 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=468970 $D=8
M1359 24041 23886 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=390500 $Y=112830 $D=8
M1360 23822 23824 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=179690 $D=8
M1361 24572 24573 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=180970 $D=8
M1362 24596 24597 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=323690 $D=8
M1363 24620 24621 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=324970 $D=8
M1364 24644 24645 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=467690 $D=8
M1365 23854 23856 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=468970 $D=8
M1366 24673 23887 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=393025 $Y=112830 $D=8
M1367 24025 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=393380 $Y=160970 $D=8
M1368 24026 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=393380 $Y=164845 $D=8
M1369 VDD 23818 23820 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=179690 $D=8
M1370 VDD 24570 24571 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=180970 $D=8
M1371 VDD 24594 24595 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=323690 $D=8
M1372 VDD 24618 24619 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=324970 $D=8
M1373 VDD 24642 24643 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=467690 $D=8
M1374 VDD 23850 23852 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=468970 $D=8
M1375 23818 23820 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=179690 $D=8
M1376 24570 24571 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=180970 $D=8
M1377 24594 24595 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=323690 $D=8
M1378 24618 24619 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=324970 $D=8
M1379 24642 24643 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=467690 $D=8
M1380 23850 23852 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=468970 $D=8
M1381 24024 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=396475 $Y=160970 $D=8
M1382 24023 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=396475 $Y=164845 $D=8
M1383 VDD 23814 23816 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=179690 $D=8
M1384 VDD 24568 24569 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=180970 $D=8
M1385 VDD 24592 24593 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=323690 $D=8
M1386 VDD 24616 24617 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=324970 $D=8
M1387 VDD 24640 24641 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=467690 $D=8
M1388 VDD 23846 23848 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=468970 $D=8
M1389 24672 23888 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=396690 $Y=112830 $D=8
M1390 23814 23816 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=179690 $D=8
M1391 24568 24569 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=180970 $D=8
M1392 24592 24593 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=323690 $D=8
M1393 24616 24617 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=324970 $D=8
M1394 24640 24641 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=467690 $D=8
M1395 23846 23848 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=468970 $D=8
M1396 24671 23889 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=399220 $Y=112830 $D=8
M1397 24021 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=399575 $Y=160970 $D=8
M1398 24022 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=399575 $Y=164845 $D=8
M1399 VDD 23810 23812 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=179690 $D=8
M1400 VDD 24566 24567 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=180970 $D=8
M1401 VDD 24590 24591 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=323690 $D=8
M1402 VDD 24614 24615 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=324970 $D=8
M1403 VDD 24638 24639 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=467690 $D=8
M1404 VDD 23842 23844 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=468970 $D=8
M1405 23810 23812 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=179690 $D=8
M1406 24566 24567 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=180970 $D=8
M1407 24590 24591 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=323690 $D=8
M1408 24614 24615 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=324970 $D=8
M1409 24638 24639 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=467690 $D=8
M1410 23842 23844 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=468970 $D=8
M1411 VDD 23806 23808 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=179690 $D=8
M1412 VDD 24564 24565 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=180970 $D=8
M1413 VDD 24588 24589 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=323690 $D=8
M1414 VDD 24612 24613 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=324970 $D=8
M1415 VDD 24636 24637 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=467690 $D=8
M1416 VDD 23838 23840 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=468970 $D=8
M1417 24020 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=402665 $Y=160970 $D=8
M1418 24019 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=402665 $Y=164845 $D=8
M1419 24670 23890 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=402880 $Y=112830 $D=8
M1420 23806 23808 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=179690 $D=8
M1421 24564 24565 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=180970 $D=8
M1422 24588 24589 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=323690 $D=8
M1423 24612 24613 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=324970 $D=8
M1424 24636 24637 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=467690 $D=8
M1425 23838 23840 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=468970 $D=8
M1426 24669 23891 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=405410 $Y=112830 $D=8
M1427 VDD 23802 23804 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=179690 $D=8
M1428 VDD 24562 24563 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=180970 $D=8
M1429 VDD 24586 24587 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=323690 $D=8
M1430 VDD 24610 24611 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=324970 $D=8
M1431 VDD 24634 24635 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=467690 $D=8
M1432 VDD 23834 23836 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=468970 $D=8
M1433 24017 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=405765 $Y=160970 $D=8
M1434 24018 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=405765 $Y=164845 $D=8
M1435 23802 23804 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=179690 $D=8
M1436 24562 24563 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=180970 $D=8
M1437 24586 24587 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=323690 $D=8
M1438 24610 24611 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=324970 $D=8
M1439 24634 24635 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=467690 $D=8
M1440 23834 23836 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=468970 $D=8
M1441 VDD 23798 23800 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=179690 $D=8
M1442 VDD 24560 24561 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=180970 $D=8
M1443 VDD 24584 24585 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=323690 $D=8
M1444 VDD 24608 24609 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=324970 $D=8
M1445 VDD 24632 24633 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=467690 $D=8
M1446 VDD 23830 23832 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=468970 $D=8
M1447 24016 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=408860 $Y=160970 $D=8
M1448 24015 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=408860 $Y=164845 $D=8
M1449 24668 23892 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=409075 $Y=112830 $D=8
M1450 23798 23800 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=179690 $D=8
M1451 24560 24561 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=180970 $D=8
M1452 24584 24585 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=323690 $D=8
M1453 24608 24609 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=324970 $D=8
M1454 24632 24633 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=467690 $D=8
M1455 23830 23832 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=468970 $D=8
M1456 VDD 23794 23796 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=179690 $D=8
M1457 VDD 24558 24559 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=180970 $D=8
M1458 VDD 24582 24583 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=323690 $D=8
M1459 VDD 24606 24607 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=324970 $D=8
M1460 VDD 24630 24631 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=467690 $D=8
M1461 VDD 23826 23828 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=468970 $D=8
M1462 24667 23893 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=411605 $Y=112830 $D=8
M1463 24013 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=411960 $Y=160970 $D=8
M1464 24014 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=411960 $Y=164845 $D=8
M1465 23794 23796 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=179690 $D=8
M1466 24558 24559 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=180970 $D=8
M1467 24582 24583 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=323690 $D=8
M1468 24606 24607 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=324970 $D=8
M1469 24630 24631 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=467690 $D=8
M1470 23826 23828 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=468970 $D=8
M1471 VDD VSS VDD VDD pfet_05v0 L=2.365e-06 W=8.19e-05 AD=0 AS=6.1309e-11 PD=0 PS=0.000217698 NRD=0 NRS=11.8457 m=1 nf=36 $X=304360 $Y=171065 $D=8
M1472 VDD VDD 23859 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=418720 $Y=467690 $D=8
M1473 VDD VDD 23857 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=418720 $Y=468970 $D=8
M1474 614 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=6.35965e-12 PD=7.86e-06 PS=1.737e-05 NRD=0.152493 NRS=0.546921 m=1 nf=2 $X=418655 $Y=160970 $D=8
M1475 615 1062 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=6.35965e-12 PD=7.86e-06 PS=1.737e-05 NRD=0.152493 NRS=0.546921 m=1 nf=2 $X=418655 $Y=164845 $D=8
M1476 23860 VSS VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=419860 $Y=467690 $D=8
M1477 23858 VSS VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=419860 $Y=468970 $D=8
M1478 606 614 VDD VDD pfet_05v0 L=6e-07 W=7.02e-06 AD=1.8252e-12 AS=3.0888e-12 PD=8.06e-06 PS=1.58e-05 NRD=0.148148 NRS=0.250712 m=1 nf=2 $X=418770 $Y=97440 $D=8
M1479 607 606 VDD VDD pfet_05v0 L=6e-07 W=2.128e-05 AD=5.5328e-12 AS=9.3632e-12 PD=2.232e-05 PS=4.432e-05 NRD=0.0488722 NRS=0.0827068 m=1 nf=2 $X=418790 $Y=67070 $D=8
M1480 613 VDD VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=2.33887e-12 PD=4.29e-06 PS=9.09e-06 NRD=0.444444 NRS=1.06061 m=1 nf=2 $X=418870 $Y=112830 $D=8
X1488 614 614 613 VDD pfet_05v0_I13 $T=419815 124190 0 180 $X=418175 $Y=116760
X1489 615 615 613 VDD pfet_05v0_I13 $T=419815 151940 0 180 $X=418175 $Y=144510
X1490 615 614 1062 VDD pfet_05v0_I13 $T=419825 159875 0 180 $X=418185 $Y=152445
X1491 614 614 VDD VSS nfet_05v0_I02 $T=419815 133465 0 180 $X=418535 $Y=126035
X1492 615 615 VDD VSS nfet_05v0_I02 $T=419815 143485 0 180 $X=418535 $Y=136055
X1498 VDD 618 616 pmos_1p2$$46273580 $T=242390 65835 1 0 $X=240960 $Y=64015
X1499 VSS 617 1000 VSS nmos_1p2$$46563372 $T=233925 66830 0 0 $X=232780 $Y=66145
X1500 618 VSS 616 VSS nmos_1p2$$46563372 $T=243510 68190 1 0 $X=242365 $Y=66555
X1501 619 618 617 VSS nmos_1p2$$46563372 $T=246080 68190 1 0 $X=244935 $Y=66555
X1503 1063 VSS Q[0] D[0] 23198 1 VDD 1064 1065 WEN[0] 23915 23916 23917 23918 23919 23920 23921 23922 23923 23924
+ 23925 23926 23927 23928 24034 1053 23885 23884 23883 23882 23881 23880 23879 23878 23877 24138 24139 24140 24141 24142
+ 24143 24144
+ saout_m2 $T=9775 25090 0 0 $X=8430 $Y=7315
X1504 1032 VSS Q[2] D[2] 23199 1 VDD 1066 1067 WEN[2] 23929 23930 23931 23932 23933 23934 23935 23936 23937 23938
+ 23939 23940 23941 23942 24035 1053 23885 23884 23883 23882 23881 23880 23879 23878 23877 24145 24146 24147 24148 24149
+ 24150 24151
+ saout_m2 $T=63775 25090 0 0 $X=62430 $Y=7315
X1505 1068 VSS Q[4] D[4] 23200 1 VDD 1069 1070 WEN[4] 23943 23944 23945 23946 23947 23948 23949 23950 23951 23952
+ 23953 23954 23955 23956 24036 1053 23886 23887 23888 23889 23890 23891 23892 23893 23877 24152 24153 24154 24155 24156
+ 24157 24158
+ saout_m2 $T=307655 25090 0 0 $X=306310 $Y=7315
X1506 1071 VSS Q[6] D[6] 23201 1 VDD 1072 1073 WEN[6] 23957 23958 23959 23960 23961 23962 23963 23964 23965 23966
+ 23967 23968 23969 23970 24037 1053 23886 23887 23888 23889 23890 23891 23892 23893 23877 24159 24160 24161 24162 24163
+ 24164 24165
+ saout_m2 $T=361655 25090 0 0 $X=360310 $Y=7315
X1507 VSS VSS 23337 23338 23339 23340 23341 23342 23343 23344 ICV_7 $T=27210 176130 1 180 $X=23870 $Y=175790
X1508 VSS VSS 23345 23346 23347 23348 23349 23350 23351 23352 ICV_7 $T=33210 176130 1 180 $X=29870 $Y=175790
X1509 VSS VSS 23353 23354 23355 23356 23357 23358 23359 23360 ICV_7 $T=81210 176130 1 180 $X=77870 $Y=175790
X1510 VSS VSS 23361 23362 23363 23364 23365 23366 23367 23368 ICV_7 $T=87210 176130 1 180 $X=83870 $Y=175790
X1511 VSS VSS 23369 23370 23371 23372 23373 23374 23375 23376 ICV_7 $T=325090 176130 1 180 $X=321750 $Y=175790
X1512 VSS VSS 23377 23378 23379 23380 23381 23382 23383 23384 ICV_7 $T=331090 176130 1 180 $X=327750 $Y=175790
X1513 VSS VSS 23385 23386 23387 23388 23389 23390 23391 23392 ICV_7 $T=379090 176130 1 180 $X=375750 $Y=175790
X1514 VSS VSS 23393 23394 23395 23396 23397 23398 23399 23400 ICV_7 $T=385090 176130 1 180 $X=381750 $Y=175790
X1515 VSS 1002 23401 23402 23403 23404 23405 23406 23407 23408 23409 23410 23411 23412 23413 23414 23415 23416 ICV_8 $T=313090 473130 0 180 $X=309750 $Y=468290
X1516 VSS 1002 23417 23418 23419 23420 23421 23422 23423 23424 23425 23426 23427 23428 23429 23430 23431 23432 ICV_8 $T=325090 473130 0 180 $X=321750 $Y=468290
X1520 VSS VSS 23433 23434 23435 23436 23437 23438 23439 23440 23441 23442 23443 23444 23445 23446 23447 23448 ICV_9 $T=12210 176130 1 180 $X=8870 $Y=175790
X1521 VSS VSS 23449 23450 23451 23452 23453 23454 23455 23456 23457 23458 23459 23460 23461 23462 23463 23464 ICV_9 $T=66210 176130 1 180 $X=62870 $Y=175790
X1522 VSS VSS 23465 23466 23467 23468 23469 23470 23471 23472 23473 23474 23475 23476 23477 23478 23479 23480 ICV_9 $T=310090 176130 1 180 $X=306750 $Y=175790
X1523 VSS VSS 23481 23482 23483 23484 23485 23486 23487 23488 23489 23490 23491 23492 23493 23494 23495 23496 ICV_9 $T=364090 176130 1 180 $X=360750 $Y=175790
X1528 VDD VSS 23202 23203 23204 23205 23206 23207 23208 23209 23210 23211 23212 23213 23214 23215 23216 23217 23218 23219
+ 23220 23221 23222 23223 23224 23225 23226 23227 23228 23229 23230 23231 23232 23233 23922 23921 23920 23919 23918 23917
+ 23916 23915 24166 24167 24168 24169 24170 24171 24172 24173 24174 24175 24176 24177 24178 24179 24180 24181
+ ICV_27 $T=12210 185130 1 180 $X=8870 $Y=180290
X1529 VDD VSS 23234 23235 23236 23237 23238 23239 23240 23241 23242 23243 23244 23245 23246 23247 23248 23249 23250 23251
+ 23252 23253 23254 23255 23256 23257 23258 23259 23260 23261 23262 23263 23264 23265 23922 23921 23920 23919 23918 23917
+ 23916 23915 24182 24183 24184 24185 24186 24187 24188 24189 24190 24191 24192 24193 24194 24195 24196 24197
+ ICV_27 $T=12210 329130 1 180 $X=8870 $Y=324290
X1530 VDD VSS 23202 23203 23204 23205 23206 23207 23208 23209 23210 23211 23212 23213 23214 23215 23216 23217 23218 23219
+ 23220 23221 23222 23223 23224 23225 23226 23227 23228 23229 23230 23231 23232 23233 23936 23935 23934 23933 23932 23931
+ 23930 23929 24198 24199 24200 24201 24202 24203 24204 24205 24206 24207 24208 24209 24210 24211 24212 24213
+ ICV_27 $T=66210 185130 1 180 $X=62870 $Y=180290
X1531 VDD VSS 23234 23235 23236 23237 23238 23239 23240 23241 23242 23243 23244 23245 23246 23247 23248 23249 23250 23251
+ 23252 23253 23254 23255 23256 23257 23258 23259 23260 23261 23262 23263 23264 23265 23936 23935 23934 23933 23932 23931
+ 23930 23929 24214 24215 24216 24217 24218 24219 24220 24221 24222 24223 24224 24225 24226 24227 24228 24229
+ ICV_27 $T=66210 329130 1 180 $X=62870 $Y=324290
X1532 VDD VSS 23266 23267 23268 23269 23270 23271 23272 23273 23274 23275 23276 23277 23278 23279 23280 23281 23282 23283
+ 23284 23285 23286 23287 23288 23289 23290 23291 23292 23293 23294 23295 23296 23297 23964 23963 23962 23961 23960 23959
+ 23958 23957 24230 24231 24232 24233 24234 24235 24236 24237 24238 24239 24240 24241 24242 24243 24244 24245
+ ICV_27 $T=364090 185130 1 180 $X=360750 $Y=180290
X1533 VDD VSS 23298 23299 23300 23301 23302 23303 23304 23305 23306 23307 23308 23309 23310 23311 23312 23313 23314 23315
+ 23316 23317 23318 23319 23320 23321 23322 23323 23324 23325 23326 23327 23328 23329 23964 23963 23962 23961 23960 23959
+ 23958 23957 24246 24247 24248 24249 24250 24251 24252 24253 24254 24255 24256 24257 24258 24259 24260 24261
+ ICV_27 $T=364090 329130 1 180 $X=360750 $Y=324290
X1534 VSS VSS 23505 23506 23507 23508 23509 23510 23511 23512 23513 23514 23515 23516 23517 23518 23519 23520 23521 23522
+ 23523 23524 23525 23526 23527 23528 23529 23530 23531 23532 23533 23534 23535 23536
+ ICV_10 $T=12210 473130 0 180 $X=8870 $Y=468290
X1535 VSS VSS 23537 23538 23539 23540 23541 23542 23543 23544 23545 23546 23547 23548 23549 23550 23551 23552 23553 23554
+ 23555 23556 23557 23558 23559 23560 23561 23562 23563 23564 23565 23566 23567 23568
+ ICV_10 $T=39210 176130 1 180 $X=35870 $Y=175790
X1536 VSS VSS 23569 23570 23571 23572 23573 23574 23575 23576 23577 23578 23579 23580 23581 23582 23583 23584 23585 23586
+ 23587 23588 23589 23590 23591 23592 23593 23594 23595 23596 23597 23598 23599 23600
+ ICV_10 $T=39210 473130 0 180 $X=35870 $Y=468290
X1537 VSS VSS 23601 23602 23603 23604 23605 23606 23607 23608 23609 23610 23611 23612 23613 23614 23615 23616 23617 23618
+ 23619 23620 23621 23622 23623 23624 23625 23626 23627 23628 23629 23630 23631 23632
+ ICV_10 $T=66210 473130 0 180 $X=62870 $Y=468290
X1538 VSS VSS 23633 23634 23635 23636 23637 23638 23639 23640 23641 23642 23643 23644 23645 23646 23647 23648 23649 23650
+ 23651 23652 23653 23654 23655 23656 23657 23658 23659 23660 23661 23662 23663 23664
+ ICV_10 $T=93210 176130 1 180 $X=89870 $Y=175790
X1539 VSS VSS 23665 23666 23667 23668 23669 23670 23671 23672 23673 23674 23675 23676 23677 23678 23679 23680 23681 23682
+ 23683 23684 23685 23686 23687 23688 23689 23690 23691 23692 23693 23694 23695 23696
+ ICV_10 $T=93210 473130 0 180 $X=89870 $Y=468290
X1540 VSS VSS 23697 23698 23699 23700 23701 23702 23703 23704 23705 23706 23707 23708 23709 23710 23711 23712 23713 23714
+ 23715 23716 23717 23718 23719 23720 23721 23722 23723 23724 23725 23726 23727 23728
+ ICV_10 $T=337090 176130 1 180 $X=333750 $Y=175790
X1541 VSS 1002 23729 23730 23731 23732 23733 23734 23735 23736 23737 23738 23739 23740 23741 23742 23743 23744 23745 23746
+ 23747 23748 23749 23750 23751 23752 23753 23754 23755 23756 23757 23758 23759 23760
+ ICV_10 $T=337090 473130 0 180 $X=333750 $Y=468290
X1542 VSS 1002 23761 23762 23763 23764 23765 23766 23767 23768 23769 23770 23771 23772 23773 23774 23775 23776 23777 23778
+ 23779 23780 23781 23782 23783 23784 23785 23786 23787 23788 23789 23790 23791 23792
+ ICV_10 $T=364090 473130 0 180 $X=360750 $Y=468290
X1543 VSS VSS 23793 23794 23795 23796 23797 23798 23799 23800 23801 23802 23803 23804 23805 23806 23807 23808 23809 23810
+ 23811 23812 23813 23814 23815 23816 23817 23818 23819 23820 23821 23822 23823 23824
+ ICV_10 $T=391090 176130 1 180 $X=387750 $Y=175790
X1544 VSS 1002 23825 23826 23827 23828 23829 23830 23831 23832 23833 23834 23835 23836 23837 23838 23839 23840 23841 23842
+ 23843 23844 23845 23846 23847 23848 23849 23850 23851 23852 23853 23854 23855 23856
+ ICV_10 $T=391090 473130 0 180 $X=387750 $Y=468290
X1568 VDD VSS 23202 23203 23204 23205 23206 23207 23208 23209 23210 23211 23212 23213 23214 23215 23216 23217 23218 23219
+ 23220 23221 23222 23223 23224 23225 23226 23227 23228 23229 23230 23231 23232 23233 23923 23924 23925 23926 23927 23928
+ 1065 1064 1076 1077 23984 23983 23982 23981 23980 23979 23978 23977 23976 23975 23974 23973 23972 23971 24262 24263
+ 24264 24265 24266 24267 24268 24269 24270 24271 24272 24273 24274 24275 24276 24277 24278 24279 24280 24281 24282 24283
+ 24284 24285 24286 24287 24288 24289 24290 24291 24292 24293 24294 24295 24296 24297 24298 24299 24300 24301 24302 24303
+ 24304 24305 24306 24307 24308 24309
+ ICV_24 $T=24210 180630 0 0 $X=23870 $Y=180290
X1569 VDD VSS 23234 23235 23236 23237 23238 23239 23240 23241 23242 23243 23244 23245 23246 23247 23248 23249 23250 23251
+ 23252 23253 23254 23255 23256 23257 23258 23259 23260 23261 23262 23263 23264 23265 23923 23924 23925 23926 23927 23928
+ 1065 1064 1076 1077 23984 23983 23982 23981 23980 23979 23978 23977 23976 23975 23974 23973 23972 23971 24310 24311
+ 24312 24313 24314 24315 24316 24317 24318 24319 24320 24321 24322 24323 24324 24325 24326 24327 24328 24329 24330 24331
+ 24332 24333 24334 24335 24336 24337 24338 24339 24340 24341 24342 24343 24344 24345 24346 24347 24348 24349 24350 24351
+ 24352 24353 24354 24355 24356 24357
+ ICV_24 $T=24210 324630 0 0 $X=23870 $Y=324290
X1570 VDD VSS 23202 23203 23204 23205 23206 23207 23208 23209 23210 23211 23212 23213 23214 23215 23216 23217 23218 23219
+ 23220 23221 23222 23223 23224 23225 23226 23227 23228 23229 23230 23231 23232 23233 23937 23938 23939 23940 23941 23942
+ 1067 1066 1079 1080 23998 23997 23996 23995 23994 23993 23992 23991 23990 23989 23988 23987 23986 23985 24358 24359
+ 24360 24361 24362 24363 24364 24365 24366 24367 24368 24369 24370 24371 24372 24373 24374 24375 24376 24377 24378 24379
+ 24380 24381 24382 24383 24384 24385 24386 24387 24388 24389 24390 24391 24392 24393 24394 24395 24396 24397 24398 24399
+ 24400 24401 24402 24403 24404 24405
+ ICV_24 $T=78210 180630 0 0 $X=77870 $Y=180290
X1571 VDD VSS 23234 23235 23236 23237 23238 23239 23240 23241 23242 23243 23244 23245 23246 23247 23248 23249 23250 23251
+ 23252 23253 23254 23255 23256 23257 23258 23259 23260 23261 23262 23263 23264 23265 23937 23938 23939 23940 23941 23942
+ 1067 1066 1079 1080 23998 23997 23996 23995 23994 23993 23992 23991 23990 23989 23988 23987 23986 23985 24406 24407
+ 24408 24409 24410 24411 24412 24413 24414 24415 24416 24417 24418 24419 24420 24421 24422 24423 24424 24425 24426 24427
+ 24428 24429 24430 24431 24432 24433 24434 24435 24436 24437 24438 24439 24440 24441 24442 24443 24444 24445 24446 24447
+ 24448 24449 24450 24451 24452 24453
+ ICV_24 $T=78210 324630 0 0 $X=77870 $Y=324290
X1572 VDD VSS 23266 23267 23268 23269 23270 23271 23272 23273 23274 23275 23276 23277 23278 23279 23280 23281 23282 23283
+ 23284 23285 23286 23287 23288 23289 23290 23291 23292 23293 23294 23295 23296 23297 23951 23952 23953 23954 23955 23956
+ 1070 1069 1083 1084 24012 24011 24010 24009 24008 24007 24006 24005 24004 24003 24002 24001 24000 23999 24454 24455
+ 24456 24457 24458 24459 24460 24461 24462 24463 24464 24465 24466 24467 24468 24469 24470 24471 24472 24473 24474 24475
+ 24476 24477 24478 24479 24480 24481 24482 24483 24484 24485 24486 24487 24488 24489 24490 24491 24492 24493 24494 24495
+ 24496 24497 24498 24499 24500 24501
+ ICV_24 $T=322090 180630 0 0 $X=321750 $Y=180290
X1573 VDD VSS 23298 23299 23300 23301 23302 23303 23304 23305 23306 23307 23308 23309 23310 23311 23312 23313 23314 23315
+ 23316 23317 23318 23319 23320 23321 23322 23323 23324 23325 23326 23327 23328 23329 23951 23952 23953 23954 23955 23956
+ 1070 1069 1083 1084 24012 24011 24010 24009 24008 24007 24006 24005 24004 24003 24002 24001 24000 23999 24502 24503
+ 24504 24505 24506 24507 24508 24509 24510 24511 24512 24513 24514 24515 24516 24517 24518 24519 24520 24521 24522 24523
+ 24524 24525 24526 24527 24528 24529 24530 24531 24532 24533 24534 24535 24536 24537 24538 24539 24540 24541 24542 24543
+ 24544 24545 24546 24547 24548 24549
+ ICV_24 $T=322090 324630 0 0 $X=321750 $Y=324290
X1574 VDD VSS 23266 23267 23268 23269 23270 23271 23272 23273 23274 23275 23276 23277 23278 23279 23280 23281 23282 23283
+ 23284 23285 23286 23287 23288 23289 23290 23291 23292 23293 23294 23295 23296 23297 23965 23966 23967 23968 23969 23970
+ 1073 1072 1086 1087 24026 24025 24024 24023 24022 24021 24020 24019 24018 24017 24016 24015 24014 24013 24550 24551
+ 24552 24553 24554 24555 24556 24557 24558 24559 24560 24561 24562 24563 24564 24565 24566 24567 24568 24569 24570 24571
+ 24572 24573 24574 24575 24576 24577 24578 24579 24580 24581 24582 24583 24584 24585 24586 24587 24588 24589 24590 24591
+ 24592 24593 24594 24595 24596 24597
+ ICV_24 $T=376090 180630 0 0 $X=375750 $Y=180290
X1575 VDD VSS 23298 23299 23300 23301 23302 23303 23304 23305 23306 23307 23308 23309 23310 23311 23312 23313 23314 23315
+ 23316 23317 23318 23319 23320 23321 23322 23323 23324 23325 23326 23327 23328 23329 23965 23966 23967 23968 23969 23970
+ 1073 1072 1086 1087 24026 24025 24024 24023 24022 24021 24020 24019 24018 24017 24016 24015 24014 24013 24598 24599
+ 24600 24601 24602 24603 24604 24605 24606 24607 24608 24609 24610 24611 24612 24613 24614 24615 24616 24617 24618 24619
+ 24620 24621 24622 24623 24624 24625 24626 24627 24628 24629 24630 24631 24632 24633 24634 24635 24636 24637 24638 24639
+ 24640 24641 24642 24643 24644 24645
+ ICV_24 $T=376090 324630 0 0 $X=375750 $Y=324290
X1576 1075 VSS Q[1] 1074 D[1] 1 VDD 1076 1077 WEN[1] 23971 23972 23973 23974 23975 23976 23977 23978 23979 23980
+ 23981 23982 23983 23984 24038 1053 23878 23879 23880 23881 23882 23883 23884 23885 23877 24646 24647 24648 24649 24650
+ 24651 24652
+ saout_R_m2 $T=65645 25125 1 180 $X=27480 $Y=6815
X1577 1033 VSS Q[3] 1078 D[3] 1 VDD 1079 1080 WEN[3] 23985 23986 23987 23988 23989 23990 23991 23992 23993 23994
+ 23995 23996 23997 23998 24039 1053 23878 23879 23880 23881 23882 23883 23884 23885 23877 24653 24654 24655 24656 24657
+ 24658 24659
+ saout_R_m2 $T=119645 25125 1 180 $X=81480 $Y=6815
X1578 1082 VSS Q[5] 1081 D[5] 1 VDD 1083 1084 WEN[5] 23999 24000 24001 24002 24003 24004 24005 24006 24007 24008
+ 24009 24010 24011 24012 24040 1053 23893 23892 23891 23890 23889 23888 23887 23886 23877 24660 24661 24662 24663 24664
+ 24665 24666
+ saout_R_m2 $T=363525 25125 1 180 $X=325360 $Y=6815
X1579 1085 VSS Q[7] 1062 D[7] 1 VDD 1086 1087 WEN[7] 24013 24014 24015 24016 24017 24018 24019 24020 24021 24022
+ 24023 24024 24025 24026 24041 1053 23893 23892 23891 23890 23889 23888 23887 23886 23877 24667 24668 24669 24670 24671
+ 24672 24673
+ saout_R_m2 $T=417525 25125 1 180 $X=379360 $Y=6815
X1581 VDD VSS 702 703 24674 24675 24676 24677 ICV_41 $T=117210 185130 0 0 $X=116870 $Y=180290
X1582 VDD VSS 702 703 24678 24679 24680 24681 ICV_41 $T=117210 221130 0 0 $X=116870 $Y=216290
X1583 VDD VSS 702 703 24682 24683 24684 24685 ICV_41 $T=117210 257130 0 0 $X=116870 $Y=252290
X1584 VDD VSS 702 703 24686 24687 24688 24689 ICV_41 $T=117210 293130 0 0 $X=116870 $Y=288290
X1585 VDD VSS 702 703 24690 24691 24692 24693 ICV_41 $T=117210 329130 0 0 $X=116870 $Y=324290
X1586 VDD VSS 702 703 24694 24695 24696 24697 ICV_41 $T=117210 365130 0 0 $X=116870 $Y=360290
X1587 VDD VSS 702 703 24698 24699 24700 24701 ICV_41 $T=117210 401130 0 0 $X=116870 $Y=396290
X1588 VDD VSS 702 703 24702 24703 24704 24705 ICV_41 $T=117210 437130 0 0 $X=116870 $Y=432290
X1589 VSS VDD 1040 1044 1046 1047 1048 1049 1050 1051 23203 23204 23205 23206 23207 23208 23267 23268 23269 23270
+ 23271 23272 1 24042 24043 24044 24045 24106 24107 24108 24109
+ ICV_37 $T=154400 190385 1 270 $X=126565 $Y=179495
X1590 VSS VDD 1040 1043 1046 1047 1048 1049 1050 1051 23211 23212 23213 23214 23215 23216 23275 23276 23277 23278
+ 23279 23280 1 24046 24047 24048 24049 24110 24111 24112 24113
+ ICV_37 $T=154400 226385 1 270 $X=126565 $Y=215495
X1591 VSS VDD 1040 1042 1046 1047 1048 1049 1050 1051 23219 23220 23221 23222 23223 23224 23283 23284 23285 23286
+ 23287 23288 1 24050 24051 24052 24053 24114 24115 24116 24117
+ ICV_37 $T=154400 262385 1 270 $X=126565 $Y=251495
X1592 VSS VDD 1040 1041 1046 1047 1048 1049 1050 1051 23227 23228 23229 23230 23231 23232 23291 23292 23293 23294
+ 23295 23296 1 24054 24055 24056 24057 24118 24119 24120 24121
+ ICV_37 $T=154400 298385 1 270 $X=126565 $Y=287495
X1593 VSS VDD 1038 1044 1046 1047 1048 1049 1050 1051 23235 23236 23237 23238 23239 23240 23299 23300 23301 23302
+ 23303 23304 1 24058 24059 24060 24061 24122 24123 24124 24125
+ ICV_37 $T=154400 334385 1 270 $X=126565 $Y=323495
X1594 VSS VDD 1038 1043 1046 1047 1048 1049 1050 1051 23243 23244 23245 23246 23247 23248 23307 23308 23309 23310
+ 23311 23312 1 24062 24063 24064 24065 24126 24127 24128 24129
+ ICV_37 $T=154400 370385 1 270 $X=126565 $Y=359495
X1595 VSS VDD 1038 1042 1046 1047 1048 1049 1050 1051 23251 23252 23253 23254 23255 23256 23315 23316 23317 23318
+ 23319 23320 1 24066 24067 24068 24069 24130 24131 24132 24133
+ ICV_37 $T=154400 406385 1 270 $X=126565 $Y=395495
X1596 VSS VDD 1038 1041 1046 1047 1048 1049 1050 1051 23259 23260 23261 23262 23263 23264 23323 23324 23325 23326
+ 23327 23328 1 24070 24071 24072 24073 24134 24135 24136 24137
+ ICV_37 $T=154400 442385 1 270 $X=126565 $Y=431495
X1600 VSS VDD 1 CLK VSS A[8] 23902 23903 1038 1040 xpredec0 $T=146075 111460 0 0 $X=144630 $Y=111455
X1601 VSS VDD 1 CLK A[7] A[6] 1041 1042 1043 1044 xpredec0 $T=182970 111460 0 0 $X=181525 $Y=111455
X1606 VSS VDD 1 CLK 23884 23885 23878 23879 23880 23881 23882 23883 23893 23892 23891 23890 23889 23888 23887 23886
+ A[2] A[1] A[0]
+ ypredec1 $T=145470 26355 0 0 $X=146365 $Y=26735
X1609 1001 VSS 1003 nfet_05v0_I20 $T=175115 470995 0 90 $X=164385 $Y=470315
X1610 1002 VSS 1004 nfet_05v0_I20 $T=260115 470995 0 90 $X=249385 $Y=470315
X1614 VDD 1001 1003 pmos_1p2_02_R90 $T=189610 471150 0 90 $X=176320 $Y=469670
X1615 VDD 1002 1004 pmos_1p2_02_R90 $T=248135 471150 0 90 $X=234845 $Y=469670
X1616 1003 VDD 2 VDD pfet_05v0_I14 $T=198405 470995 0 90 $X=191195 $Y=469955
X1617 1 2 VSS VDD pfet_05v0_I14 $T=219905 470995 0 90 $X=212695 $Y=469955
X1618 1004 VDD 2 VDD pfet_05v0_I14 $T=233255 470995 0 90 $X=226045 $Y=469955
X1619 1003 VSS 2 nfet_05v0_I11 $T=202950 470995 0 90 $X=199690 $Y=470315
X1620 1004 VSS 2 nfet_05v0_I11 $T=224800 470995 0 90 $X=221540 $Y=470315
X1621 VSS VDD GWEN CLK 23877 1053 wen_v2 $T=208415 16605 0 0 $X=208280 $Y=15275
X1622 VSS 1 VDD CLK A[5] A[4] A[3] 1045 1046 1047 1048 1049 1050 1051 1052 xpredec1 $T=219860 111460 0 0 $X=219855 $Y=111455
X1623 VDD 1005 CLK pfet_05v0_I08 $T=234280 43425 1 0 $X=233240 $Y=41905
X1624 VDD 1006 1005 pfet_05v0_I08 $T=239670 43425 1 0 $X=238630 $Y=41905
X1625 VSS 1005 CLK nfet_05v0_I15 $T=234280 46585 1 0 $X=233600 $Y=45365
X1626 VSS 1006 1005 nfet_05v0_I15 $T=239670 46585 1 0 $X=238990 $Y=45365
X1638 VDD VSS 23266 23267 23268 23269 23270 23271 23272 23273 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24738 24739 24740 24741 24742 24743 24744 24745 24746 24747 24748 24749 24750 24751 24752 24753 24754 24755 24756 24757
+ ICV_31 $T=307090 180630 1 180 $X=303750 $Y=180290
X1639 VDD VSS 23274 23275 23276 23277 23278 23279 23280 23281 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24758 24759 24760 24761 24762 24763 24764 24765 24766 24767 24768 24769 24770 24771 24772 24773 24774 24775 24776 24777
+ ICV_31 $T=307090 216630 1 180 $X=303750 $Y=216290
X1640 VDD VSS 23282 23283 23284 23285 23286 23287 23288 23289 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24778 24779 24780 24781 24782 24783 24784 24785 24786 24787 24788 24789 24790 24791 24792 24793 24794 24795 24796 24797
+ ICV_31 $T=307090 252630 1 180 $X=303750 $Y=252290
X1641 VDD VSS 23290 23291 23292 23293 23294 23295 23296 23297 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24798 24799 24800 24801 24802 24803 24804 24805 24806 24807 24808 24809 24810 24811 24812 24813 24814 24815 24816 24817
+ ICV_31 $T=307090 288630 1 180 $X=303750 $Y=288290
X1642 VDD VSS 23298 23299 23300 23301 23302 23303 23304 23305 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24818 24819 24820 24821 24822 24823 24824 24825 24826 24827 24828 24829 24830 24831 24832 24833 24834 24835 24836 24837
+ ICV_31 $T=307090 324630 1 180 $X=303750 $Y=324290
X1643 VDD VSS 23306 23307 23308 23309 23310 23311 23312 23313 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24838 24839 24840 24841 24842 24843 24844 24845 24846 24847 24848 24849 24850 24851 24852 24853 24854 24855 24856 24857
+ ICV_31 $T=307090 360630 1 180 $X=303750 $Y=360290
X1644 VDD VSS 23314 23315 23316 23317 23318 23319 23320 23321 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24858 24859 24860 24861 24862 24863 24864 24865 24866 24867 24868 24869 24870 24871 24872 24873 24874 24875 24876 24877
+ ICV_31 $T=307090 396630 1 180 $X=303750 $Y=396290
X1645 VDD VSS 23322 23323 23324 23325 23326 23327 23328 23329 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24878 24879 24880 24881 24882 24883 24884 24885 24886 24887 24888 24889 24890 24891 24892 24893 24894 24895 24896 24897
+ ICV_31 $T=307090 432630 1 180 $X=303750 $Y=432290
X1648 614 615 VSS VDD 24074 24075 24076 24077 ICV_4 $T=415090 176130 0 0 $X=414750 $Y=175790
X1649 614 615 VSS VDD 24078 24079 24080 24081 ICV_4 $T=415090 212130 0 0 $X=414750 $Y=211790
X1650 614 615 VSS VDD 24082 24083 24084 24085 ICV_4 $T=415090 248130 0 0 $X=414750 $Y=247790
X1651 614 615 VSS VDD 24086 24087 24088 24089 ICV_4 $T=415090 284130 0 0 $X=414750 $Y=283790
X1652 614 615 VSS VDD 24090 24091 24092 24093 ICV_4 $T=415090 320130 0 0 $X=414750 $Y=319790
X1653 614 615 VSS VDD 24094 24095 24096 24097 ICV_4 $T=415090 356130 0 0 $X=414750 $Y=355790
X1654 614 615 VSS VDD 24098 24099 24100 24101 ICV_4 $T=415090 392130 0 0 $X=414750 $Y=391790
X1655 614 615 VSS VDD 24102 24103 24104 24105 ICV_4 $T=415090 428130 0 0 $X=414750 $Y=427790
.ENDS
