* Subcircuit definition of cell ICV_26
.SUBCKT ICV_26 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 36 37 38 39 40 41 42 43 44 45 46 47 48 49
+ 50 51
** N=67 EP=42 IP=80 FDC=368
*.SEEDPROM
M0 7 58 59 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-11370 $Y=30560 $D=8
M1 7 66 67 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-11370 $Y=31840 $D=8
M2 58 59 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-10230 $Y=30560 $D=8
M3 66 67 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-10230 $Y=31840 $D=8
M4 7 56 57 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=30560 $D=8
M5 7 64 65 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=31840 $D=8
M6 56 57 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=30560 $D=8
M7 64 65 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=31840 $D=8
M8 7 54 55 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=30560 $D=8
M9 7 62 63 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=31840 $D=8
M10 54 55 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=30560 $D=8
M11 62 63 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=31840 $D=8
M12 7 52 53 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=30560 $D=8
M13 7 60 61 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=31840 $D=8
M14 52 53 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=30560 $D=8
M15 60 61 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=31840 $D=8
X16 7 8 9 10 11 12 13 14 15 16 32 31 30 29 28 27 26 25 36 37
+ 38 39 40 41 42 43 52 53 54 55 56 57 58 59
+ ICV_25 $T=0 0 0 0 $X=-12340 $Y=-4840
X17 7 8 17 18 19 20 21 22 23 24 32 31 30 29 28 27 26 25 60 61
+ 62 63 64 65 66 67 44 45 46 47 48 49 50 51
+ ICV_25 $T=0 36000 0 0 $X=-12340 $Y=31160
.ENDS
