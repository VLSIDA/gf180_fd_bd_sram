* Subcircuit definition of cell pmoscap_L1_W2_R270
.SUBCKT pmoscap_L1_W2_R270
** N=13 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
