* Subcircuit definition of cell xdec32
.SUBCKT xdec32 vss xc xb[3] xb[2] xb[1] xb[0] xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] xa[1] xa[0] vdd LWL[0] LWL[1] LWL[2] LWL[3] LWL[4]
+ LWL[5] LWL[6] LWL[7] LWL[8] LWL[9] LWL[10] LWL[11] LWL[12] LWL[13] LWL[14] LWL[15] LWL[16] LWL[17] LWL[18] LWL[19] LWL[20] LWL[21] LWL[22] LWL[23] LWL[24]
+ LWL[25] LWL[26] LWL[27] LWL[28] LWL[29] LWL[30] LWL[31] RWL[1] RWL[2] RWL[3] RWL[4] RWL[5] RWL[6] RWL[7] RWL[8] RWL[9] RWL[10] RWL[11] RWL[12] RWL[13]
+ RWL[14] RWL[15] RWL[16] RWL[17] RWL[18] RWL[19] RWL[20] RWL[21] RWL[22] RWL[23] RWL[24] RWL[25] RWL[26] RWL[27] RWL[28] RWL[29] RWL[30] RWL[31] RWL[0] men
** N=357 EP=80 IP=544 FDC=608
M0 vss 326 LWL[0] vss nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=16340 $Y=260 $D=2
M1 326 310 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=2660 $D=2
M2 vss 312 328 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=32740 $D=2
M3 vss 328 LWL[7] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=34020 $D=2
M4 vss 330 LWL[8] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=36260 $D=2
M5 330 314 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=38660 $D=2
M6 vss 316 332 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=68740 $D=2
M7 vss 332 LWL[15] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=70020 $D=2
M8 vss 334 LWL[16] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=72260 $D=2
M9 334 318 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=74660 $D=2
M10 vss 320 336 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=104740 $D=2
M11 vss 336 LWL[23] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=106020 $D=2
M12 vss 338 LWL[24] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=108260 $D=2
M13 338 322 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=110660 $D=2
M14 vss 324 340 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=140740 $D=2
M15 vss 340 LWL[31] vss nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=16340 $Y=142020 $D=2
M16 310 311 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=46620 $Y=260 $D=2
M17 vss 313 312 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=46620 $Y=35140 $D=2
M18 314 315 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=46620 $Y=36260 $D=2
M19 vss 317 316 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=46620 $Y=71140 $D=2
M20 318 319 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=46620 $Y=72260 $D=2
M21 vss 321 320 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=46620 $Y=107140 $D=2
M22 322 323 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=46620 $Y=108260 $D=2
M23 vss 325 324 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=46620 $Y=143140 $D=2
M24 343 xc vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=7.32375e-13 AS=2.079e-12 PD=3.615e-06 PS=7.62e-06 NRD=0.0738095 NRS=0.209524 m=1 nf=1 $X=66460 $Y=315 $D=2
M25 342 xb[0] 343 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=1380 $D=2
M26 311 xa[0] 342 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=2500 $D=2
M27 344 xa[7] 313 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=32900 $D=2
M28 345 xb[0] 344 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=34020 $D=2
M29 vss xc 345 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=66460 $Y=35085 $D=2
M30 347 xc vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=66460 $Y=36315 $D=2
M31 346 xb[1] 347 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=37380 $D=2
M32 315 xa[0] 346 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=38500 $D=2
M33 348 xa[7] 317 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=68900 $D=2
M34 349 xb[1] 348 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=70020 $D=2
M35 vss xc 349 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=66460 $Y=71085 $D=2
M36 351 xc vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=66460 $Y=72315 $D=2
M37 350 xb[2] 351 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=73380 $D=2
M38 319 xa[0] 350 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=74500 $D=2
M39 352 xa[7] 321 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=104900 $D=2
M40 353 xb[2] 352 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=106020 $D=2
M41 vss xc 353 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=66460 $Y=107085 $D=2
M42 355 xc vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=66460 $Y=108315 $D=2
M43 354 xb[3] 355 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=109380 $D=2
M44 323 xa[0] 354 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=110500 $D=2
M45 356 xa[7] 325 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=140900 $D=2
M46 357 xb[3] 356 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=142020 $D=2
M47 vss xc 357 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.079e-12 AS=7.32375e-13 PD=7.62e-06 PS=3.615e-06 NRD=0.209524 NRS=0.0738095 m=1 nf=1 $X=66460 $Y=143085 $D=2
M48 vss 327 RWL[0] vss nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=100255 $Y=260 $D=2
M49 327 310 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=2660 $D=2
M50 vss 312 329 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=32740 $D=2
M51 vss 329 RWL[7] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=34020 $D=2
M52 vss 331 RWL[8] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=36260 $D=2
M53 331 314 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=38660 $D=2
M54 vss 316 333 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=68740 $D=2
M55 vss 333 RWL[15] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=70020 $D=2
M56 vss 335 RWL[16] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=72260 $D=2
M57 335 318 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=74660 $D=2
M58 vss 320 337 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=104740 $D=2
M59 vss 337 RWL[23] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=106020 $D=2
M60 vss 339 RWL[24] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=108260 $D=2
M61 339 322 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=110660 $D=2
M62 vss 324 341 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=140740 $D=2
M63 vss 341 RWL[31] vss nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=100255 $Y=142020 $D=2
M64 vdd 326 LWL[0] vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=4665 $Y=260 $D=8
M65 LWL[7] 328 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=4665 $Y=32900 $D=8
M66 vdd 330 LWL[8] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=4665 $Y=36260 $D=8
M67 LWL[15] 332 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=4665 $Y=68900 $D=8
M68 vdd 334 LWL[16] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=4665 $Y=72260 $D=8
M69 LWL[23] 336 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=4665 $Y=104900 $D=8
M70 vdd 338 LWL[24] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=4665 $Y=108260 $D=8
M71 LWL[31] 340 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=4665 $Y=140900 $D=8
M72 311 xc vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=260 $D=8
M73 vdd xb[0] 311 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=1380 $D=8
M74 311 xa[0] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=2500 $D=8
M75 vdd xa[7] 313 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=32900 $D=8
M76 313 xb[0] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=34020 $D=8
M77 vdd xc 313 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=35140 $D=8
M78 315 xc vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=36260 $D=8
M79 vdd xb[1] 315 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=37380 $D=8
M80 315 xa[0] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=38500 $D=8
M81 vdd xa[7] 317 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=68900 $D=8
M82 317 xb[1] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=70020 $D=8
M83 vdd xc 317 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=71140 $D=8
M84 319 xc vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=72260 $D=8
M85 vdd xb[2] 319 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=73380 $D=8
M86 319 xa[0] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=74500 $D=8
M87 vdd xa[7] 321 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=104900 $D=8
M88 321 xb[2] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=106020 $D=8
M89 vdd xc 321 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=107140 $D=8
M90 323 xc vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=108260 $D=8
M91 vdd xb[3] 323 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=109380 $D=8
M92 323 xa[0] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=110500 $D=8
M93 vdd xa[7] 325 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=140900 $D=8
M94 325 xb[3] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=142020 $D=8
M95 vdd xc 325 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=143140 $D=8
M96 vdd 327 RWL[0] vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=106930 $Y=260 $D=8
M97 RWL[7] 329 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=106930 $Y=32900 $D=8
M98 vdd 331 RWL[8] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=106930 $Y=36260 $D=8
M99 RWL[15] 333 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=106930 $Y=68900 $D=8
M100 vdd 335 RWL[16] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=106930 $Y=72260 $D=8
M101 RWL[23] 337 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=106930 $Y=104900 $D=8
M102 vdd 339 RWL[24] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=106930 $Y=108260 $D=8
M103 RWL[31] 341 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=106930 $Y=140900 $D=8
X104 vss xc xb[0] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] vdd 310 men 311 LWL[1] RWL[1] LWL[2] RWL[2] LWL[3] RWL[3] LWL[4]
+ RWL[4] LWL[5] RWL[5] LWL[6] RWL[6] 312 313 326 327 328 329
+ xdec8 $T=0 0 0 0 $X=0 $Y=-1140
X105 vss xc xb[1] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] vdd 314 men 315 LWL[9] RWL[9] LWL[10] RWL[10] LWL[11] RWL[11] LWL[12]
+ RWL[12] LWL[13] RWL[13] LWL[14] RWL[14] 316 317 330 331 332 333
+ xdec8 $T=0 36000 0 0 $X=0 $Y=34860
X106 vss xc xb[2] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] vdd 318 men 319 LWL[17] RWL[17] LWL[18] RWL[18] LWL[19] RWL[19] LWL[20]
+ RWL[20] LWL[21] RWL[21] LWL[22] RWL[22] 320 321 334 335 336 337
+ xdec8 $T=0 72000 0 0 $X=0 $Y=70860
X107 vss xc xb[3] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] vdd 322 men 323 LWL[25] RWL[25] LWL[26] RWL[26] LWL[27] RWL[27] LWL[28]
+ RWL[28] LWL[29] RWL[29] LWL[30] RWL[30] 324 325 338 339 340 341
+ xdec8 $T=0 108000 0 0 $X=0 $Y=106860
.ENDS
