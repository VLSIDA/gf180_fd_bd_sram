* Subcircuit definition of cell pfet_05v0_I10
.SUBCKT pfet_05v0_I10
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
