* Subcircuit definition of cell ICV_11
.SUBCKT ICV_11
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
