* Subcircuit definition of cell pmos_1p2$$202587180
.SUBCKT pmos_1p2$$202587180
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
