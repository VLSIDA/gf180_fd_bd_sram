* Subcircuit definition of cell ICV_7
.SUBCKT ICV_7 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
** N=30 EP=18 IP=33 FDC=16
*.SEEDPROM
X0 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 ICV_5 $T=-3000 0 0 0 $X=-12340 $Y=-340
.ENDS
