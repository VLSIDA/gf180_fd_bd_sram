* Subcircuit definition of cell ICV_20
.SUBCKT ICV_20
** N=6 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
