* Subcircuit definition of cell ICV_35
.SUBCKT ICV_35 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32
+ 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52
+ 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72
+ 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92
+ 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112
+ 113 114 115 116 117 118
** N=118 EP=106 IP=168 FDC=704
*.SEEDPROM
X0 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 55 56
+ 57 58 59 60 61 62 63 64 65 66 67 68 69 70
+ ICV_34 $T=-42000 -4500 0 0 $X=-51340 $Y=-4840
X1 13 14 15 16 17 18 19 20 21 22 31 32 33 34 35 36 37 38 71 72
+ 73 74 75 76 77 78 79 80 81 82 83 84 85 86
+ ICV_34 $T=-30000 -4500 0 0 $X=-39340 $Y=-4840
X4 13 14 15 16 17 18 19 20 21 22 39 40 41 42 43 44 45 46 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ ICV_30 $T=-12000 -4500 1 180 $X=-24340 $Y=-4840
X5 13 14 15 16 17 18 19 20 21 22 47 48 49 50 51 52 53 54 103 104
+ 105 106 107 108 109 110 111 112 113 114 115 116 117 118
+ ICV_30 $T=0 -4500 1 180 $X=-12340 $Y=-4840
.ENDS
