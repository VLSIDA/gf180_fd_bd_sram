* Subcircuit definition of cell ICV_16
.SUBCKT ICV_16
** N=15 EP=0 IP=20 FDC=0
.ENDS
