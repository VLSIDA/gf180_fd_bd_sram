* Subcircuit definition of cell xpredec0
.SUBCKT xpredec0 vss vdd men clk A[1] A[0] x[3] x[2] x[1] x[0]
** N=99 EP=10 IP=158 FDC=56
M0 x[3] 90 vss vss nfet_05v0 L=6e-07 W=1.816e-05 AD=4.7216e-12 AS=5.5388e-12 PD=2.024e-05 PS=2.514e-05 NRD=0.229075 NRS=0.268722 m=1 nf=4 $X=260 $Y=50820 $D=2
M1 x[2] 92 vss vss nfet_05v0 L=6e-07 W=1.816e-05 AD=4.7216e-12 AS=4.7216e-12 PD=2.024e-05 PS=2.024e-05 NRD=0.229075 NRS=0.229075 m=1 nf=4 $X=4740 $Y=50820 $D=2
M2 x[1] 94 vss vss nfet_05v0 L=6e-07 W=1.816e-05 AD=4.7216e-12 AS=4.7216e-12 PD=2.024e-05 PS=2.024e-05 NRD=0.229075 NRS=0.229075 m=1 nf=4 $X=9220 $Y=50820 $D=2
M3 x[0] 96 vss vss nfet_05v0 L=6e-07 W=1.816e-05 AD=4.7216e-12 AS=5.5388e-12 PD=2.024e-05 PS=2.514e-05 NRD=0.229075 NRS=0.268722 m=1 nf=4 $X=13700 $Y=50820 $D=2
M4 17 men vss vss nfet_05v0 L=6e-07 W=1.37e-06 AD=3.562e-13 AS=6.028e-13 PD=1.89e-06 PS=3.62e-06 NRD=0.189781 NRS=0.321168 m=1 nf=1 $X=21630 $Y=51200 $D=2
M5 vss clk 17 vss nfet_05v0 L=6e-07 W=1.37e-06 AD=6.028e-13 AS=3.562e-13 PD=3.62e-06 PS=1.89e-06 NRD=0.321168 NRS=0.189781 m=1 nf=1 $X=22750 $Y=51200 $D=2
M6 x[3] 90 vdd vdd pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.38348e-11 PD=4.744e-05 PS=5.914e-05 NRD=0.0917108 NRS=0.107584 m=1 nf=4 $X=260 $Y=38080 $D=8
M7 x[2] 92 vdd vdd pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.744e-05 PS=4.744e-05 NRD=0.0917108 NRS=0.0917108 m=1 nf=4 $X=4740 $Y=38080 $D=8
M8 x[1] 94 vdd vdd pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.744e-05 PS=4.744e-05 NRD=0.0917108 NRS=0.0917108 m=1 nf=4 $X=9220 $Y=38080 $D=8
M9 x[0] 96 vdd vdd pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.38348e-11 PD=4.744e-05 PS=5.914e-05 NRD=0.0917108 NRS=0.107584 m=1 nf=4 $X=13700 $Y=38080 $D=8
M10 98 men vdd vdd pfet_05v0 L=6e-07 W=1.705e-06 AD=4.39037e-13 AS=1.01447e-12 PD=2.22e-06 PS=4.6e-06 NRD=0.151026 NRS=0.348974 m=1 nf=1 $X=21630 $Y=47525 $D=8
M11 17 clk 98 vdd pfet_05v0 L=6e-07 W=1.705e-06 AD=8.525e-15 AS=-8.525e-15 PD=1e-08 PS=-1e-08 NRD=0.00293255 NRS=-0.00293255 m=1 nf=1 $X=22745 $Y=47525 $D=8
M12 99 clk 17 vdd pfet_05v0 L=6e-07 W=1.705e-06 AD=-8.525e-15 AS=8.525e-15 PD=-1e-08 PS=1e-08 NRD=-0.00293255 NRS=0.00293255 m=1 nf=1 $X=23870 $Y=47525 $D=8
M13 vdd men 99 vdd pfet_05v0 L=6e-07 W=1.705e-06 AD=1.01447e-12 AS=4.39037e-13 PD=4.6e-06 PS=2.22e-06 NRD=0.348974 NRS=0.151026 m=1 nf=1 $X=24985 $Y=47525 $D=8
M14 18 17 vdd vdd pfet_05v0 L=6e-07 W=2.28e-06 AD=5.928e-13 AS=1.0032e-12 PD=3.32e-06 PS=6.32e-06 NRD=0.45614 NRS=0.77193 m=1 nf=2 $X=29010 $Y=47595 $D=8
X17 18 vss 17 vss nmos_1p2$$46563372 $T=29755 51180 0 0 $X=28610 $Y=50495
X18 90 vss vdd 30 31 xpredec0_xa $T=-2205 170 0 0 $X=-1440 $Y=-5
X19 92 vss vdd 30 32 xpredec0_xa $T=11165 170 1 180 $X=3000 $Y=-5
X20 94 vss vdd 33 31 xpredec0_xa $T=6755 170 0 0 $X=7520 $Y=-5
X21 96 vss vdd 33 32 xpredec0_xa $T=20125 170 1 180 $X=11960 $Y=-5
X22 vss 30 33 vdd A[1] 17 18 xpredec0_bot $T=18665 3160 0 0 $X=18135 $Y=-5
X23 vss 31 32 vdd A[0] 17 18 xpredec0_bot $T=27120 3160 0 0 $X=26590 $Y=-5
.ENDS
