* Subcircuit definition of cell pmos_1p2$$47815724
.SUBCKT pmos_1p2$$47815724
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
