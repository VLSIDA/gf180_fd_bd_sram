* Subcircuit definition of cell M1_PSUB$$47122476
.SUBCKT M1_PSUB$$47122476
** N=5 EP=0 IP=0 FDC=0
.ENDS
