* Subcircuit definition of cell din
.SUBCKT din vss 2 3 4 5 6 7 8 d db 11 12 vdd datain men wep
** N=69 EP=16 IP=73 FDC=24
M0 2 4 vss vss nfet_05v0 L=6e-07 W=1.361e-05 AD=5.9884e-12 AS=5.9884e-12 PD=2.81e-05 PS=2.81e-05 NRD=0.0323292 NRS=0.0323292 m=1 nf=1 $X=260 $Y=10430 $D=2
M1 3 wep vss vss nfet_05v0 L=6e-07 W=1.14e-06 AD=7.866e-13 AS=7.923e-13 PD=3.66e-06 PS=3.67e-06 NRD=0.605263 NRS=0.609649 m=1 nf=1 $X=3600 $Y=38320 $D=2
M2 vss 7 4 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=11165 $Y=8655 $D=2
M3 3 wep vdd vdd pfet_05v0 L=6e-07 W=2.97e-06 AD=1.13602e-12 AS=1.7523e-12 PD=4.5e-06 PS=8.3e-06 NRD=0.515152 NRS=0.794613 m=1 nf=2 $X=3025 $Y=35440 $D=8
M4 vdd 2 11 vdd pfet_05v0 L=6e-07 W=1.134e-05 AD=4.9896e-12 AS=4.9896e-12 PD=2.356e-05 PS=2.356e-05 NRD=0.0388007 NRS=0.0388007 m=1 nf=1 $X=6980 $Y=26220 $D=8
X5 4 vdd 7 vdd pfet_05v0_I01 $T=11165 455 0 0 $X=10125 $Y=-165
X6 d 2 3 vdd pmos_1p2$$46889004 $T=2655 26220 0 0 $X=1225 $Y=25510
X7 db 11 3 vdd pmos_1p2$$46889004 $T=4895 26220 0 0 $X=3465 $Y=25510
X10 5 vss 6 datain 5 vss nfet_05v0_I11 $T=2765 1790 1 0 $X=2085 $Y=210
X11 6 7 8 12 men vss nfet_05v0_I11 $T=6905 725 0 0 $X=6225 $Y=105
X12 d 2 wep vss nmos_1p2$$46883884 $T=2655 12695 0 0 $X=1510 $Y=12010
X13 db 11 wep vss nmos_1p2$$46883884 $T=4895 12695 0 0 $X=3750 $Y=12010
X14 11 vss 2 vss nmos_1p2$$46883884 $T=7135 12695 0 0 $X=5990 $Y=12010
X15 vss 12 men vss nmos_1p2$$46563372 $T=3470 9035 0 0 $X=2325 $Y=8350
X16 vss 8 4 vss nmos_1p2$$46563372 $T=7060 10495 1 0 $X=5915 $Y=8860
X17 5 vdd 6 datain 5 vdd pfet_05v0_I18 $T=2765 3195 0 0 $X=1725 $Y=2575
X18 6 7 8 men 12 vdd pfet_05v0_I18 $T=6905 3605 0 0 $X=5865 $Y=2985
X19 vdd 12 men pmos_1p2$$46273580 $T=2920 7175 1 0 $X=1490 $Y=5355
X20 vdd 8 4 pmos_1p2$$46273580 $T=7060 8140 1 0 $X=5630 $Y=6320
X21 vdd 2 4 pmos_1p2$$46887980 $T=415 26220 0 0 $X=-1015 $Y=25510
.ENDS
