* Subcircuit definition of cell ypredec1_bot
.SUBCKT ypredec1_bot 1 2 3 10 11 12 13
** N=34 EP=7 IP=20 FDC=12
M0 2 30 1 1 nfet_05v0 L=6e-07 W=4.54e-06 AD=1.9976e-12 AS=1.9976e-12 PD=9.96e-06 PS=9.96e-06 NRD=0.0969163 NRS=0.0969163 m=1 nf=1 $X=3755 $Y=33350 $D=2
M1 3 2 1 1 nfet_05v0 L=6e-07 W=4.54e-06 AD=1.9976e-12 AS=1.9976e-12 PD=9.96e-06 PS=9.96e-06 NRD=0.0969163 NRS=0.0969163 m=1 nf=1 $X=6325 $Y=33350 $D=2
X2 10 2 30 pmos_1p2$$46887980 $T=3910 18340 0 0 $X=2480 $Y=17630
X3 10 3 2 pmos_1p2$$46887980 $T=6480 18340 0 0 $X=5050 $Y=17630
X6 1 30 11 10 13 12 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
.ENDS
